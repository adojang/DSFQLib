.title KiCad schematic
R3 /11x /10a Resistor
RB1 /10a /102 Resistor
L1 A /10 Inductor
LJ1 /101 /3 Inductor
B1 /101 /10a jjmit
PLR1 /100 /3 Inductor
R1 /10 /100 Resistor
LCa1 /10 /10a Inductor
LC1 /3 /7 Inductor
PRB1 /102 /3 Inductor
LC5 /7 /8 Inductor
LJ5 /80 /90 Inductor
B5 /80 /8 jjmit
PRB5 /81 /90 Inductor
RB5 /8 /81 Resistor
L3 /8 Q Inductor
LRBias1 Bias /8 Resistor
LP1 /90 GND Inductor
RB4 /21 /221 Resistor
PRB4 /221 /7 Inductor
LJ3 /110 /7 Inductor
LJ4 /220 /7 Inductor
PLR3 /11x /11 Inductor
B3 /110 /11 jjmit
B4 /220 /21 jjmit
PLR4 /21x /21 Inductor
PRB3 /111 /7 Inductor
RB3 /11 /111 Resistor
R4 /21x /20a Resistor
PRB2 /202 /5 Inductor
LC2 /5 /7 Inductor
B2 /201 /20a jjmit
RB2 /20a /202 Resistor
LJ2 /201 /5 Inductor
PLR2 /200 /5 Inductor
R2 /20 /200 Resistor
L2 B /20 Inductor
LCb1 /20 /20a Inductor
.end
