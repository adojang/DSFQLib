* DSFQ Self clocked Multiplexor
* Author: Adriaan van Wijk
* Version: 1.0
* Last modification date: 21 June 2022
* Last modification by: Adriaan van Wijk
* This testbench uses cells from LS's library of RSFQ cells. This was the version that was tested for layout.

.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include cells\AW_mitll_OR_optimized.cir
.include cells\AW_mitll_AND_optimized.cir
.include cells\LSmitll_SPLIT_v2p1_optimized.cir
.include cells\LSmitll_NOT_v2p1_optimized.cir


.param cval=600u


I_a0 0 I_a0 pwl(0 0 200p 0 203p cval 205p 0 300p 0 303p cval 305p 0)
I_b0 0 I_b0 pwl(0 0 85p 0 88p cval 90p 0 300p 0 303p cval 305p 0)
*IMPORTANT! The s0 line requires VERY fine timing for the NOT gate to work. It might be worth adding something on both ends of the NOT gate to enable a little bit of play. It will extend the time the not gate takes to trigger, but it will probably be worth it.

I_s0 0 I_s0 pwl(0 0 107p 0 110p cval 112p 0 307p 0 310p cval 312p 0)
*S = 0 - Select A
*S = 1 - Select B

*I_s0 0 I_s0 pwl(0 0 200p 0 203p cval 205p 0 300p 0 303p cval 305p 0)


.tran 0.25p 1500p 0 0.01p

Xsrc_a0 LSmitll_DCSFQ i_a0 src_a0
Xsrc_b0 LSmitll_DCSFQ i_b0 src_b0
Xsrc_s0 LSmitll_DCSFQ i_s0 src_s0

Xload_a0 LSMITLL_JTL src_a0 A0
Xload_b0 LSMITLL_JTL src_b0 B0
Xload_s0 LSMITLL_JTL src_s0 S0

XSPLITA LSMITLL_SPLIT A0 A1 A_clk
XSPLITB LSMITLL_SPLIT B0 B1 B_clk
XSPLITS LSMITLL_SPLIT S0 S1 B2

XORCLK  DSFQ_OR    A_clk B_clk CLK
XCLKBOOST LSMITLL_JTL CLK CLK_BOOST

XNOT    LSMITLL_NOT   S1 CLK_BOOST A2

XAND1   DSFQ_AND   A1 A2 Q1
XAND2   DSFQ_AND   B1 B2 Q2

XOR     DSFQ_OR    Q1 Q2 QQ


Xloadout_s0 LSMITLL_JTL QQ Qload
R_out Qload 0 2



.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)


*.print v(A0) v(B0) v(S1) v(CLK) v(A2) v(S0) v(R_out)
.print v(A1) v(S1) v(CLK_BOOST) v(A2) p(Q1) p(Q2) p(QQ)
.end