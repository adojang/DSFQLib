.title KiCad schematic
L4 /5 /9 Inductor
I1 GND /9 pwl(0 0 5p REF)
L3 CLK /5 Inductor
L5 /9 /10 Inductor
LP1 /6 GND Inductor
B5 /6 /5 jjmit
L6 /10 /11 Inductor
L2 A /4 Inductor
B4 /12 /11 jjmit
B6 /7 /10 jjmit
LP2 /7 GND Inductor
L7 /12 /13 Inductor
B3 /12 /4 jjmit
L10 /17 Q Inductor
L8 /13 /16 Inductor
LP5 /8 GND Inductor
B9 /8 /12 jjmit
I3 GND /4 pwl(0 0 5p REF)
L9 /16 /17 Inductor
I2 GND /16 pwl(0 0 5p REF)
LP4 /15 GND Inductor
B8 /15 /17 jjmit
B7 /14 /13 jjmit
LP3 /14 GND Inductor
.end
