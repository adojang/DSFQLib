*25.8% Skew for a tolerance of 15ps
.subckt DSFQ_OR a b q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

*Confluence Buffer A

.param l1   =     1.64019283e-12
.param b1   =     2.40525670e+00
.param b3   =     2.98576249e+00
.param b4   =     4.08935660e-01


* AND GATE LOOP
.param l4   =     1.08922491e-12
.param b7   =     1.47293130e+00
.param b9   =     5.33372490e-01
.param lr2   =     1.48265019e-13
.param r1   =     5.59076275e+00
.param r2   =     4.90609696e-01
.param lr1   =     5.08374673e-13


* Output Stage
.param b8   =     4.27449779e-01
.param i1   =     3.07565196e-04
.param l3   =     1.79574511e-12
.param l6   =     2.00183654e-12


*Confluence Buffer B
.param 	l2  	= L1
.param 	b2  	= B1
.param 	b5  	= B3
.param 	b6  	= B4

*Parasitics
.param 	lp1  	= 0.2e-12
.param 	lp2  	= 0.2e-12
.param 	lp3  	= 0.2e-12
.param 	lp5  	= 0.2e-12

* Back Annotated .cir file from KiCad
b1   	1   	1j   	 jjmit area=b1
b2   	2   	2j   	 jjmit area=b2
b3   	10   	3   	 jjmit area=b3
b4   	3   	5   	 jjmit area=b4
b5   	10   	4   	 jjmit area=b5
b6   	4   	6   	 jjmit area=b6
b7   	20   	24   	 jjmit area=b7
b8   	30   	31   	 jjmit area=b8
b9   	23   	24   	 jjmit area=b9

i1   	0   	10   	pwl(0   	0   	5p      i1)
l1   	a   	1   	 l1
l2   	b   	2   	 l2
l3   	10   	30   	 l3
l4   	30   	20   	 l4
l6   	30   	q   	 l6

LJ1     1j      3       0
LJ2     2j      4       0

lR1   	21   	24   	 lr1
lR2   	22   	23   	 LR2


lp1   	5   	0   	 lp1
lp2   	6   	0   	 lp2
lp3   	24   	0   	 lp3
lp5   	31   	0   	 lp5
r1   	21   	20   	 r1
r2   	22   	20   	 r2
.ends