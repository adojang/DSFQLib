* JSIM deck file generated with TimEx
* === DEVICE-UNDER-TEST ===

* === SOURCE DEFINITION ===
.SUBCKT SOURCECELL  8 11
b1   1  2  jjmitll100 area=2.25
b2   3  4  jjmitll100 area=2.25
b3   5  6  jjmitll100 area=2.5
ib1  0  2  pwl(0 0 5p 275ua)
ib2  0  5  pwl(0 0 5p 175ua)
l1   8  7  1p
l2   7  0  3.9p
l3   7  1  0.6p
l4   2  3  1.1p
l5   3  5  4.5p
l6   5  11 2p
lp2  4  0  0.2p
lp3  6  0  0.2p
lrb1 9  2  1p
lrb2 10 4  1p
lrb3 12 6  1p
rb1  1  9  4.31
rb2  3  10 4.31
rb3  5  12 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS SOURCECELL
* === INPUT LOAD DEFINITION ===
.SUBCKT LOADINCELL  2 5
b1 1 6 jjmitll100 area=2.5
b2 4 8 jjmitll100 area=2.5
ib1 0 3 pwl(0 0 5p 350ua)
l1 2 1 2p
l2 1 3 2p
l3 3 4 2p
l4 4 5 2p
lb1 7 6 1p
lb2 9 8 1p
lp1 6 0 0.2p
lp2 8 0 0.2p
rb1 1 7 3.88
rb2 4 9 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS LOADINCELL
* === OUTPUT LOAD DEFINITION ===
.SUBCKT LOADOUTCELL  2 5
b1 1 6 jjmitll100 area=2.5
b2 4 8 jjmitll100 area=2.5
ib1 0 3 pwl(0 0 5p 350ua)
l1 2 1 2p
l2 1 3 2p
l3 3 4 2p
l4 4 5 2p
lb1 7 6 1p
lb2 9 8 1p
lp1 6 0 0.2p
lp2 8 0 0.2p
rb1 1 7 3.88
rb2 4 9 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS LOADOUTCELL
* === SINK DEFINITION ===
.SUBCKT SINKCELL  1
r1 1 0 2
.ENDS SINKCELL
* ===== MAIN =====
.param cval=600u
I_a 0 1000 pwl(0 0 
+100p 0 103p cval 105p 0 
+400p 0 403p cval 405p 0
+500p 0 503p cval 505p 0
+515p 0 518p cval 520p 0
+615p 0 618p cval 620p 0
+860p 0 863p cval 865p 0)

I_b 0 4000 pulse(cval 0 200p 1p 1p 3p 200p)

.tran 0.25p 1000p 0 0.01p

XSOURCEINa SOURCECELL 1000 2000
XLOADINa LOADINCELL 2000 A

XSOURCEINb SOURCECELL 4000 5000
XLOADINb LOADINCELL 5000 B
XLOADOUTq LOADOUTCELL q 8000
XSINKOUTq SINKCELL 8000

*Optimized OR Gate

XDUT DSFQ_OR A B q

*$Ports 		 A B q
.subckt DSFQ_OR A B q

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)


*There is not enough current flowing through Blb to trigger it. LBias must increase.
.param B_JIA=    1.08172342e+00
.param B_JUA=    9.98731934e-01
.param B_JLA=    9.61678975e-01

.param B_JIB=    9.77749297e-01
.param B_JUB=    1.09557322e+00
.param B_JLB=    1.16185870e+00 

.param B_JP =    5.19248148e-01
.param B_JPS =   4.07603769e-01
.param B_JLIM=   1.96555868e+00 

.param Ibias=    2.53670849e-04 

.param LBias=    3.46560565e-10
.param Lpoff=    1.29760632e-11
.param Rs   =    9.90210690e-01 
.param RH   =    2.95746005e+00 

.param LP  =     8.19946788e-13
.param RP  =     1.08687967e+00


B_JIA A 1   jjmit area=B_JIA
B_JUA 1 N   jjmit area=B_JUA
B_JLA 1 0   jjmit area=B_JLA

B_JIB B 3   jjmit area=B_JIB
B_JUB 3 N   jjmit area=B_JUB
B_JLB 3 0   jjmit area=B_JLB

B_JP 4 0    jjmit area=B_JP
B_JPS 5 0   jjmit area=B_JPS

B_JLIM 2 6  jjmit area=B_JLIM

Lpoff 2 4 Lpoff
Rs 4 5 Rs
RH 4 0 RH

Lbias 0 6 Lbias
Lcon N 2 4p
IBM 0 N pwl(0 0 5p Ibias)

*Parasitic Inductances and Resistances for each JJ
RJIA A 1a RP
RJUA 1 Na RP
RJLA 1 G1 RP

RJIB B 3b RP
RJUB 3 Nb RP
RJLB 3 G3 RP

RJP 4 G4 RP
RJPS 5 G5 RP

RJLIM 2 6q RP

LJIA 1a 1   LP
LJUA Na N   LP
LJLA G1 0   LP

LJIB 3b 3   LP
LJUB Nb N   LP
LJLB G3 0   LP

LJP  G4 0   LP
LJPS G5 0   LP

LJLIM 6q 6  LP

Lout 2 q 2p
.ends


.print v(L4.XLOADINa) v(L4.XLOADINb) v(Lout.XDUT) p(r1.XSINKOUTq)
.end
