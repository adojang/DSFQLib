.include LSmitll_MERGE_v2p1_optimized.cir
.include LSmitll_XOR_v2p1_optimized.cir
.include LSmitll_SPLIT_v2p1_optimized.cir

*Propagation Delay Times:
*XSPLIT -   12ps
*XMRG   -   9ps
*XOR    -   16ps
*Total =    28ps (longest path XSPLIT-XOR)

.subckt DSFQ_XOR A B q


XSPLITA LSmitll_SPLIT A A1 A2
XSPLITB LSmitll_SPLIT B B1 B2
XMRGCLK LSmitll_MERGE A2 B2 MRGCLK
XXOR LSmitll_XOR A1 B1 MRGCLK q
.ends