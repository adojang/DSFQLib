.title KiCad schematic
B5 /31 /30 jjmit
RB5 /30 /32 Resistor
LP1 /31 GND Inductor
LRB5 /32 GND Inductor
R4 /22 /20 Resistor
R1 /10 /30 Resistor
B1 /30 /10 jjmit
B3 /30 /12 jjmit
B2 /30 /20 jjmit
B4 /30 /22 jjmit
R2 /20 /30 Resistor
L1 A /10 Inductor
R3 /12 /10 Resistor
L2 B /20 Inductor
L3 /30 /40 Inductor
I1 GND /30 pwl(0 0 5p REF)
B7 /41 /40 jjmit
LRB7 /42 GND Inductor
LP7 /41 GND Inductor
L4 /50 /51 Inductor
RB6 /50 /43 Resistor
RB7 /40 /42 Resistor
B6 /40 /50 jjmit
LRB6 /43 /40 Inductor
L5 /40 D Inductor
L6 /51 C Inductor
I2 GND /51 pwl(0 0 5p REF)
.end
