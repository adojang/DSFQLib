* A Generic Testbench for simulating Logic Gates
* Copyright (c) 2022-2024 Adriaan van Wijk, Stellenbosch University
*
*
* This testbench is not meant to be attached to PTLs as it does not support integrated PTL ports.
*
*
*
*
*


*===== SFQ Source =======
*$Ports 			a q
.subckt LSmitll_DCSFQ a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

.param B0=1.0
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LB=2p
.param LP=0.2p

.param B1=2.25
.param B2=2.25
.param B3=2.5
.param L1=1p
.param L2=3.9p
.param L3=0.6p
.param L4=1.1p
.param L5=4.5p
.param L6=2p
.param IB1=275u
.param IB2=175u
.param LB1=LB
.param LB2=LB
.param LP2=LP
.param LP3=LP
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet

B1 2 3 jjmit area=B1
B2 5 6 jjmit area=B2
B3 7 8 jjmit area=B3
IB1 0 4 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
LB1 3 4 LB1
LB2 7 9 LB2
L1 a 1 L1
L2 1 0 L2
L3 1 2 L3
L4 3 5 L4
L5 5 7 L5
L6 7 q L6
LP2 6 0 LP2
LP3 8 0 LP3
RB1 2 102 RB1
LRB1 102 3 LRB1
RB2 5 105 RB2
LRB2 105 0 LRB2
RB3 7 107 RB3
LRB3 107 0 LRB3

.ends

*=========== JTL LOADS ==========
*$Ports 			a q
.subckt LSMITLL_JTL a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=IC
.param IB1=(B1+B2)*Ic0*BiasCoef
.param LB1=LB
.param L1=Phi0/(4*B1*Ic0)
.param L2=Phi0/(4*B1*Ic0)
.param L3=Phi0/(4*B1*Ic0)
.param L4=Phi0/(4*B2*Ic0)
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP

B1 1 2 jjmit area=B1
B2 6 7 jjmit area=B2
IB1 0 5 pwl(0 0 5p IB1)
L1 a 1 L1
L2 1 4 L2
L3 4 6 L3
L4 6 q L4
LP1 2 0 LP1
LP2 7 0 LP2
LB1 5 4 LB1
RB1 1 3 RB1
RB2 6 8 RB2
LRB1 3 0 LRB1
LRB2 8 0 LRB2

.ends

*====== Device Under Test ======
*$Ports 		 A B Q
.subckt DSFQ_AND A B Q

.model main jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=84uA)
.model secondary jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=60uA)
.model third jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=168uA)

L1 A 1 12p
L2 B 4 12p
RD1 1 2 0.67 neb=10G
RD2 4 5 0.67 neb=10G
BD1 2 C secondary
BD2 5 C secondary
B1 1 C main
B2 4 C main
B3 C 0 third

Ibias 0 C dc 70u

.ends

*=========== END DUT =========

*====== Main TestBench========


XSourceA LSmitll_DCSFQ srcAin srcAout
XSourceB LSmitll_DCSFQ srcBin srcBout

XLoadInA LSMITLL_JTL srcaout loadaout
XLoadInB LSMITLL_JTL srcbout loadbout

*=======================================
XDUT DSFQ_AND loadaout loadbout dutout
*=======================================

XLoadCircuit LSMITLL_JTL dutout loadout
RSink loadout 0 2

* ==SOURCE CURRENT INPUTS==

* The tests below are preconfigured for common logic gate tests.
* The tests include timing tests which are neccesary for DSFQ to be verified.
* If two inputs arrive within X time of one another, both are considered (nominally 40ps)

.param cval = 700u


* BASIC Timing Tests are each 100ps apart:
*IsrcA 0 srcain pwl(0 0 100p 0 101p cval 102p 0 300p 0 301p cval 302p 0)
*IsrcB 0 srcbin pwl(0 0 200p 0 201p cval 202p 0 300p 0 301p cval 302p 0)

* BASIC Timing Tests each 50ps apart:
*IsrcA 0 srcain pwl(0 0 50p 0 51p cval 52p 0 150p 0 151p cval 152p 0)
*IsrcB 0 srcbin pwl(0 0 100p 0 101p cval 102p 0 150p 0 151p cval 152p 0)

* Advanced Tests to see how long a value is held 20ps 30ps 40ps
IsrcA 0 srcain pwl(0 0 50p 0 51p cval 52p 0 150p 0 151p cval 152p 0 250p 0 251p cval 252p 0)
IsrcB 0 srcbin pwl(0 0 70p 0 71p cval 72p 0 180p 0 181p 0 182p 0 290p 0 291p cval 292p 0)

*Note that with these settings, the trigger is somehow 'held back' for an extended period. This may be a design issue.


* Advanced Tests to demonstrate multiple input rejection



.tran 0.25p 500p 0 0.01p

*Prints Circuit Inputs, and Circuit Output
.print i(L6.XSourceA) i(L6.XSourceB) i(RSink) p(B3.XDUT) p(B1.XLoadCircuit)
.end