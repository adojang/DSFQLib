* Author: Adriaan van Wijk
* Version: 1.0
* Last modification date: 21 Feburary 2021
* Last modification by: Adriaan van Wijk
* Based on the design by Rylov [2019]

* Copyright (c) 2021 Adriaan van Wijk, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Adriaan van Wijk, 21786275@sun.ac.za


*$Ports 		 A B q
.subckt DSFQ_OR A B q

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)


.param B_JIA    =   1.2
.param B_JUA    =   1
.param B_JLA    =   1.3

.param B_JIB    =   1.2
.param B_JUB    =   1
.param B_JLB    =   1.3

.param B_JP     =   0.7
.param B_PS     =   0.5
.param B_JLIM   =   1.8

.param Ibias = 250u

.param LBias    =   350p
.param Lpoff    =   16p
.param Rs=1
.param RH=4

.param LP       =   1p
.param RP       =   1


B_JIA A 1   jjmit area=B_JIA
B_JUA 1 N   jjmit area=B_JUA
B_JLA 1 0   jjmit area=B_JLA

B_JIB B 3   jjmit area=B_JIB
B_JUB 3 N   jjmit area=B_JUB
B_JLB 3 0   jjmit area=B_JLB

B_JP 4 0    jjmit area=B_JP
B_JPS 5 0   jjmit area=B_JPS

B_JLIM 2 6  jjmit area=B_JLIM

Lpoff 2 4 Lpoff
Rs 4 5 Rs
RH 4 0 RH

Lbias 0 6 Lbias
Lcon N 2 4p
IBM 0 N pwl(0 0 5p Ibias)

*Parasitic Inductances and Resistances for each JJ
RJIA A 1a RP
RJUA 1 Na RP
RJLA 1 G1 RP

RJIB B 3b RP
RJUB 3 Nb RP
RJLB 3 G3 RP

RJP 4 G4 RP
RJPS 5 G5 RP

RJLIM 2 6q RP

LJIA 1a 1   LP
LJUA Na N   LP
LJLA G1 0   LP

LJIB 3b 3   LP
LJUB Nb N   LP
LJLB G3 0   LP

LJP  G4 0   LP
LJPS G5 0   LP

LJLIM 6q 6  LP

Lout 2 q 2p
.ends