*OR Gate by Rylov.
*$Ports 		 A B q
.subckt DSFQ_OR A B q

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

.param Bps=0.5
.param Bp=0.7
.param Bia=1.2
.param Bib=1.2
.param Bua=1
.param Bub=1
.param Bla=1.3
.param Blb=1.3
.param Blim=1.8

.param LBias 350p
.param Lpoff = 16p
.param Rs=1
.param RH=4
.param IB1=270u


*Noise
*Noise
.param pinduct = 1p

Bia A 1 jjmit area=Bia
Ria A 10 1.97
Lia 10 1 pinduct

Bib B 3 jjmit area=Bib
Rib B 11 1.97
Lib 11 3 pinduct

Bua 1 2 jjmit area=Bua
Rua 1 13 2.16
Lua 13 2 pinduct

Bub 3 2 jjmit area=Bub
Rub 3 14 2.16
Lub 14 2 pinduct

Bla 1 0 jjmit area=Bla
Rla 1 15 1.90
Lla 15 0 pinduct

Blb 3 0 jjmit area=Blb
Rlb 3 16 1.90
Llb 16 0 pinduct

Lpoff 2 4 Lpoff

Rs 4 5 Rs

*Dunno if this should be here.
RH 4 0 RH

Bp 4 0 jjmit area=Bp
Rp 4 17 2.59
Lp 17 0 pinduct

Bps 5 0 jjmit area=Bps
Rps 5 18 2.79
Lps 18 0 pinduct

Lbias q VDD Lbias

*Delay of about 50ps from input to output.
*Cutoff value seems to be 260. 270 looks ideal
IB1 0 VDD (0 0 5p IB1)

Blim q 2 jjmit area=Blim
Rlim 19 2 1.6
Llim 19 q pinduct
.ends