.param 	b3  	= 1.38
.param 	b4  	= 1.36
.param 	b5  	= 1
.param 	b6  	= 1
.param 	b7  	= 1
.param 	b8  	= 1
.param 	b9  	= 0.80
.param 	i1  	= 140u
.param 	i2  	= 140u
.param 	i3  	= 100u
.param 	l10  	= 2p
.param 	l2  	= 2p
.param 	l3  	= 2p
.param 	l4  	= 2p
.param 	l5  	= 2p
.param 	l6  	= 4p
.param 	l7  	= 2p
.param 	l8  	= 2p
.param 	l9  	= 2p
.param 	lp1  	= 0.2p
.param 	lp2  	= 0.2p
.param 	lp3  	= 0.2p
.param 	lp4  	= 0.2p
.param 	lp5  	= 0.2p