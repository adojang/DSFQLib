*.subckt master a b c q
.param lad  	=	 	    5

xtest1 one a b q1
xtest2 two q1 c q

*.subckt one am bm q1m
l_connect_0 xaa xaa 0

l_connect_1 xbb xbb 0

l1 am xaa 5
r1 xbb bm 5
c1 xbb qm1
xtest3 three saa_three_one sbb_three_one


*.subckt three saa sbb
l_connect_0_three xrr_three xrr_three 0

l_connect_1_three xyy_three xyy_three 0

l1_three saa_three fr1_three 55
lr_three fr1_three xrr_three 553
lk_three xyy_three sbb_three 33

xrinox rhino oupa_rhino_three_one hannes_rhino_three_one

*.subckt rhino oupa hannes
.param opsies_rhino_three = 55
.param katjie_rhino_three = 767
r1_rhino_three oupa_rhino_three hannes_rhino_three opsies_rhino_three
r2_rhino_three hannes_rhino_three 0 katjie_rhino_three
*.ends


*.ends


*.ends

*.ends

*.ends


*.subckt two q1m cm q
l1_two q1m_two cm_two 5
r1_two q1_two 0 5
c1_two q11_two q_two *.ends_two




*.ends