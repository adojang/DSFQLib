.param 	b1  	= 
.param 	b2  	= 
.param 	b3  	= 
.param 	b4  	= 
.param 	b5  	= 
.param 	i1  	= 
.param 	l1  	= 
.param 	l2  	= 
.param 	l3  	= 
.param 	lp1  	= 
.param 	lrb1  	= 
.param 	lrb2  	= 
.param 	lrb3  	= 
.param 	lrb4  	= 
.param 	lrb5  	= 
.param 	r1  	= 
.param 	r2  	= 
.param 	r3  	= 
.param 	r4  	= 
.param 	rb1  	= 
.param 	rb2  	= 
.param 	rb3  	= 
.param 	rb4  	= 
.param 	rb5  	= 


* Back Annotated .cir file from KiCad
b1   	30   	10   	 jjmit area=b1
b2   	30   	20   	 jjmit area=b2
b3   	30   	12   	 jjmit area=b3
b4   	30   	22   	 jjmit area=b4
b5   	31   	30   	 jjmit area=b5
i1   	0   	30   	pwl(0   	0   	5p   	i1)
l1   	a   	10   	 l1
l2   	b   	20   	 l2
l3   	30   	q   	 l3
lp1   	31   	0   	 lp1
lrb1   	11   	30   	 lrb1
lrb2   	21   	30   	 lrb2
lrb3   	net-_lrb3-pad1_   	30   	 lrb3
lrb4   	net-_lrb4-pad1_   	30   	 lrb4
lrb5   	32   	0   	 lrb5
r1   	10   	30   	 r1
r2   	20   	30   	 r2
r3   	12   	10   	 r3
r4   	22   	20   	 r4
rb1   	10   	11   	 rb1
rb2   	20   	21   	 rb2
rb3   	12   	net-_lrb3-pad1_   	 rb3
rb4   	22   	net-_lrb4-pad1_   	 rb4
rb5   	30   	32   	 rb5
.end