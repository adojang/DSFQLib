* DSFQ Self clocked Multiplexor
* Author: Adriaan van Wijk
* Version: 1.0
* Last modification date: 21 June 2022
* Last modification by: Adriaan van Wijk
* This testbench uses cells from LS's library of RSFQ cells. This was the version that was tested for layout.

.include AW_mitll_DSFQ_MUX_ex.cir
.param cval=600u

I_a0 0 I_a0 pwl(0 0 100p 0 103p 0 105p 0        200p 0 203p cval 205p 0     300p 0 303p cval 305p 0     400p 0 403p 0 405p 0)
I_b0 0 I_b0 pwl(0 0 100p 0 103p cval 105p 0     200p 0 203p cval 205p 0     300p 0 303p 0 305p 0        400p 0 403p cval 405p 0)
I_s0 0 I_s0 pwl(0 0 100p 0 103p 0 105p 0        200p 0 203p 0 205p 0        300p 0 303p cval 305p 0     400p 0 403p cval 405p 0)
*S = 0 - Select A
*S = 1 - Select B

* A   0 1 1 0
* B   1 1 0 1
* S   0 0 1 1
* A2  0 1 0 0
* Q1: 0 1 0 0
* Q2: 0 0 0 1
* QQ: 0 1 0 1


.tran 0.25p 600p 0 0.01p

Xsrc_a0 LSmitll_DCSFQ i_a0 src_a0
Xsrc_b0 LSmitll_DCSFQ i_b0 src_b0
Xsrc_s0 LSmitll_DCSFQ i_s0 src_s0

Xload_a0 LSMITLL_JTL src_a0 A0
Xload_b0 LSMITLL_JTL src_b0 B0
Xload_s0 LSMITLL_JTL src_s0 S0

XMUX DSFQ_MUX A0 B0 S0 QQ
XLOAD LSMITLL_JTL QQ Qload
R_out Qload 0 2

* .print p(A0) p(B0) p(S1.xmux) p(CLK.xmux) p(B2.xmux) p(A2.xmux) p(Q1.xmux) p(Q2.xmux) p(QQ)

.print p(Q1.xmux) p(Q2.xmux) p(QQ)
