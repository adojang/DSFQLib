.include AW_mitll_AND_optimized.cir
.include AW_mitll_OR_optimized.cir
.include AW_mitll_XOR.cir
.include LSmitll_BUFF_v2p1_optimized.cir
*.include LSmitll_JTL_v2p1_optimized.cir

.subckt FULL_ADDER A B Cin Cout S
XXOR1 DSFQ_XOR A B 1
XXOR2 DSFQ_XOR 1 Cin S

XAND1 DSFQ_AND A B 3
XAND2 DSFQ_AND 1 Cin 4
XOR1 DSFQ_OR 4 3 Coutx
XSTABLE LSMITLL_JTL Coutx CoutStable
XBUFF LSMITLL_BUFF CoutStable Cout 
.ends