*DSFQ OR GATE

.model 50 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=50uA)
.model 70 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=70uA)
.model 100 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)
.model 120 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=120uA)
.model 130 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=130uA)
.model 180 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=180uA)

Bia A 1 120
Bib B 3 120
Bua 1 2 100
Bub 2 3 100
Bla 1 0 130
Blb 3 0 130

Lpoff 2 4 16p

Rs 4 5 1

Bp 4 0 70
Bps 5 0 50

Lbias 6 0 350p
Blim 2 6 180



VinA B 0 pwl(0 0 20p 0 21p 2.07m 22p 0 200p 0 201p 2.07m 202p 0)
VinB A 0 pwl(0 0 100p 0 101p 2.07m 102p 0 200p 0 201p 2.07m 202p 0)

*VDDbias vdd 0 dc 1m



.tran 0.25p 300p 0 0.01p

.print DEVI Bia
.print DEVI Bib
.print DEVI Blim
.print PHASE Blim
.end