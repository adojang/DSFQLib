.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include cells\LSmitll_SPLIT_v2p1_optimized.cir
.include cells\LSmitll_NOT_v2p1_optimized.cir
.include AW_mitll_DSFQ_AND.cir
.include AW_mitll_DSFQ_OR.cir
.include AW_mitll_DSFQ_NOT.cir
.include AW_mitll_DSFQ_XOR.cir

.param cval=600u

I_a0 0 I_a0 pwl(0 0 100p 0 103p cval 105p 0           200p 0 203p 0 205p 0         300p 0 303p cval 305p 0     400p 0 403p 0 405p 0)
I_b0 0 I_b0 pwl(0 0 100p 0 103p 0 105p 0             200p 0 203p cval 205p 0       300p 0 303p cval 305p 0     400p 0 403p 0 405p 0)

* A     0 0 1 1
* B     0 1 0 1
* AND1  0 0 0 1
* AND2  0 1 1 0
* Q     0 1 1 0


.tran 0.25p 500p 0 0.01p

Xsrc_a0 LSmitll_DCSFQ i_a0 src_a0
Xsrc_b0 LSmitll_DCSFQ i_b0 src_b0


Xload_a0 LSMITLL_JTL src_a0 A0
Xload_b0 LSMITLL_JTL src_b0 B0

XXOR DSFQ_XOR A0 B0 QQ

XLOAD LSMITLL_JTL QQ Qload
R_out Qload 0 2

.print p(A0) p(B0) p(QQ)


.end