* Author: Adriaan van Wijk
* Version: 1.4
* Last modification date: 14 April 2022
* Last modification by: Adriaan van Wijk

* Copyright (c) 2022 Adriaan van Wijk, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Adriaan van Wijk, 21786275@sun.ac.za

*********************************
* Additional Notes

* The optimized logic cell has a skew tolerance of ~ 11ps between inputs A and B.



*$Ports    A B q
.subckt DSFQ_AND A B q

.param b1       =         5.16417451e-01
.param b2       =         b1
.param b3       =         3.12658647e-01
.param b4       =         b3
.param b5       =         1.05188201e+00
.param i1       =         3.26322383e-05
.param l1       =         3.51004037e-12
.param l2       =         l1
.param l3       =         1.17410569e-12
.param lp1      =         1.40215763e-13
.param lrb1     =         2.99321337e-12
.param lrb2     =         4.83421859e-12
.param lrb3     =         3.70854087e-12
.param lrb4     =         1.79101012e-12
.param lrb5     =         1.95576828e-12
.param r1       =         1.76782953e+00
.param r2       =         r1
.param r3       =         8.40028656e-01
.param r4       =         r3
.param rb1      =         3.42859137e+00
.param rb2      =         9.41371385e+00
.param rb3      =         4.60171344e+00
.param rb4      =         5.75143516e+00
.param rb5      =         2.79007373e+00


b1   	4   	5   	 jjmit area=b1
b2   	6   	7   	 jjmit area=b2
b3   	4   	8   	 jjmit area=b3
b4   	6   	4   	 jjmit area=b4
b5   	4   	9   	 jjmit area=b5
i1   	0   	4   	pwl(0   	0   	5p   	i1)
l1   	a   	5   	 l1
l2   	b   	7   	 l2
l3   	4   	q   	 l3
lp1   	9   	0   	 lp1
lrb1   	10   	4   	 lrb1
lrb2   	11   	6   	 lrb2
lrb3   	12   	4   	 lrb3
lrb4   	13   	6   	 lrb4
lrb5   	14   	0   	 lrb5
r1   	5   	4   	 r1
r2   	7   	6   	 r2
r3   	8   	5   	 r3
r4   	4   	7   	 r4
rb1   	5   	10   	 rb1
rb2   	7   	11   	 rb2
rb3   	8   	12   	 rb3
rb4   	4   	13   	 rb4
rb5   	4   	14   	 rb5
.ends