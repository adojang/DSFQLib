* DSFQ Self clocked Multiplexor
* Author: Adriaan van Wijk
* Version: 1.0
* Last modification date: 21 June 2022
* Last modification by: Adriaan van Wijk
* This testbench uses cells from LS's library of RSFQ cells. This was the version that was tested for layout.

.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include cells\AW_mitll_OR_optimized.cir
.include cells\AW_mitll_AND_optimized.cir
.include cells\LSmitll_SPLIT_v2p1_optimized.cir
.include cells\LSmitll_NOT_v2p1_optimized.cir
.include cells\LSmitll_BUFF_v2p1_optimized.cir
.include AW_mitll_AND.cir
.include AW_mitll_INV.cir


.param cval=600u


I_a0 0 I_a0 pwl(0 0 100p 0 103p cval 105p 0 200p 0 203p cval 205p 0 300p 0 303p 0 305p 0 400p 0 403p cval 405p 0)
I_b0 0 I_b0 pwl(0 0 100p 0 103p 0 105p 0 200p 0 203p cval 205p 0 300p 0 303p cval 305p 0 400p 0 403p cval 405p 0)
I_s0 0 I_s0 pwl(0 0 100p 0 103p 0 105p 0 200p 0 203p 0 205p 0 300p 0 303p cval 305p 0 400p 0 403p cval 405p 0)
*S = 0 - Select A
*S = 1 - Select B

.tran 0.25p 500p 0 0.01p

Xsrc_a0 LSmitll_DCSFQ i_a0 src_a0
Xsrc_b0 LSmitll_DCSFQ i_b0 src_b0
Xsrc_s0 LSmitll_DCSFQ i_s0 src_s0

Xload_a0 LSMITLL_JTL src_a0 A0
Xload_b0 LSMITLL_JTL src_b0 B0
Xload_s0 LSMITLL_JTL src_s0 S0

XSPLITA LSMITLL_SPLIT A0 A1 A_clk
XSPLITB LSMITLL_SPLIT B0 B1 B_clk
XSPLITS LSMITLL_SPLIT S0 S1 B2

*XJTLQ1 LSmitll_JTL Q1 QQ1
*XJTLQ2 LSmitll_JTL Q2 QQ2

XSYNC   DSFQ_INV S1 A_clk A2

*These Shunt JJ's are required to prevent back propagation and suppress 'noise' from other signals.
B_shunts1   a_clk   	0   	 jjmit area=1.5
B_shuntQ1  	Q1   	0   	 jjmit area=1
B_shuntQ2  	Q2   	0   	 jjmit area=1
B_shuntS0   B2   	0   	 jjmit area=1.5

*Updated shuntless AND Gates 'x'
XAND1   DSFQ_ANDx   A1 A2 Q1
XAND2   DSFQ_ANDx   B1 B2 Q2

XOR     DSFQ_OR    Q1 Q2 QQ
Xloadout_s0 LSMITLL_JTL QQ Qload
R_out Qload 0 2


.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)

*.print v(A0) v(B0) v(S1) v(CLK) v(A2) v(S0) v(R_out)
*.print p(A1) p(S1) p(A_CLK) p(B1) p(B2) p(A2) p(Q1) p(Q2) p(QQ)
.print v(A0) v(B0) p(Q1) p(Q2) v(S1) p(QQ) 
*.print p(S1) p(A1) p(A2) p(a0) p(Q1) p(Q2) p(B1) p(B2)










.end