*Version Created Specifically for the DSFQ_NOT
* Hold Time of about 8ps
* Not thoroughly tested. This is a ducktape-style fix meant to be replaced later on.
.subckt DSFQ_LOOP in q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)
*8ps HOLD TIME
.param LD = 6p
.param RD = 70
.param RS = 70
LD in leak LD
RD leak d1 RD
RS leak out RS
BD d1 out jjmit area=0.7
RBD d1 gg 9.7999
LBD gg out 5.5369p
BS leak out jjmit area=1
RBS leak g9 6.8599
LBS g9 out 3.8758p
ROUT out q 0
.ends