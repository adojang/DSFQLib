.subckt DSFQ_NOT A B C Q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
*A is inverting input.
*B and C are inputs for the OR gate.
*Q is output.

XNOT LSMITLL_NOT A      CLKb    Q
XJTL LSMITLL_JTL CLKa   CLKb
XOR DSFQ_OR      B      C       CLKa

.ends
