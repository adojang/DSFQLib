.include LSmitll_MERGE_v2p1_optimized.cir
.include LSmitll_XOR_v2p1_optimized.cir
.include LSmitll_SPLIT_v2p1_optimized.cir


.subckt DSFQ_XOR A B q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)
XSPLITA LSmitll_SPLIT A A1 A2
XSPLITB LSmitll_SPLIT B B1 B2
XMRGCLK LSmitll_MERGE A2 B2 MRGCLK
XXOR LSmitll_XOR A1 B1 MRGCLK q
.ends