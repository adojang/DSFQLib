* DSFQ Self clocked Multiplexor
* Author: Adriaan van Wijk
* Version: 1.0
* Last modification date: 21 June 2022
* Last modification by: Adriaan van Wijk
* This testbench uses cells from LS's library of RSFQ cells. This was the version that was tested for layout.

.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include cells\LSmitll_SPLIT_v2p1_optimized.cir
.include cells\LSmitll_NOT_v2p1_optimized.cir
.include cells\LSmitll_BUFF_v2p1_optimized.cir
.include newadder.cir
.include AW_mitll_DSFQ_AND.cir
.include AW_mitll_DSFQ_OR.cir
.include AW_mitll_DSFQ_NOT.cir
.include AW_mitll_DSFQ_XOR.cir


.param cval=600u
I_a0 0 I_a0 pwl(0 0 200p 0 203p cval 205p 0       400p 0 403p 0 405p 0        600p 0 603p 0 605p 0        800p 0 803p cval 805p 0        1000p 0 1003p cval 1005p 0        1200p 0 1203p cval 1205p 0        1400p 0 1403p cval 1405p 0)
I_b0 0 I_b0 pwl(0 0 200p 0 203p 0 205p 0       400p 0 403p cval 405p 0        600p 0 603p cval 605p 0        800p 0 803p 0 805p 0        1000p 0 1003p 0 1005p 0        1200p 0 1203p cval 1205p 0        1400p 0 1403p cval 1405p 0)
I_ci 0 I_ci pwl(0 0 200p 0 203p cval 205p 0       400p 0 403p 0 405p 0        600p 0 603p cval 605p 0        800p 0 803p 0 805p 0        1000p 0 1003p cval 1005p 0        1200p 0 1203p 0 1205p 0        1400p 0 1403p cval 1405p 0)

I_s0 0 I_s0 pwl(0 0 200p 0 203p 0 205p 0       400p 0 403p cval 405p 0        600p 0 603p 0 605p 0        800p 0 803p cval 805p 0        1000p 0 1003p 0 1005p 0        1200p 0 1203p 0 1205p 0        1400p 0 1403p cval 1405p 0)
* I_s0 0 I_s0 pwl(0 0 170p 0 173p cval 175p 0     270p 0 273p cval 275p 0      370p 0 373p 0 375p 0        470p 0 473p cval 475p 0        570p 0 573p 0 575p 0            670p 0 673p 0 675p 0            770p 0 773p cval 775p 0)
I_z0 0 I_z0 pwl(0 0 200p 0 203p 0 205p 0       400p 0 403p 0 405p 0        600p 0 603p cval 605p 0        800p 0 803p 0 805p 0        1000p 0 1003p cval 1005p 0        1200p 0 1203p cval 1205p 0        1400p 0 1403p cval 1405p 0)



* I_a0 0 I_a0 pwl(0 0 200p 0 203p 0 205p 0       400p 0 403p 0 405p 0        600p 0 603p 0 605p 0        800p 0 803p 0 805p 0        1000p 0 1003p 0 1005p 0        1200p 0 1203p 0 1205p 0        1400p 0 1403p 0 1405p 0)
* I_b0 0 I_b0 pwl(0 0 200p 0 203p 0 205p 0       400p 0 403p 0 405p 0        600p 0 603p cval 605p 0        800p 0 803p 0 805p 0        1000p 0 1003p 0 1005p 0        1200p 0 1203p 0 1205p 0        1400p 0 1403p 0 1405p 0)
* I_ci 0 I_ci pwl(0 0 200p 0 203p 0 205p 0       400p 0 403p 0 405p 0        600p 0 603p cval 605p 0        800p 0 803p 0 805p 0        1000p 0 1003p 0 1005p 0        1200p 0 1203p 0 1205p 0        1400p 0 1403p 0 1405p 0)

* I_s0 0 I_s0 pwl(0 0 200p 0 203p cval 205p 0       400p 0 403p cval 405p 0        600p 0 603p 0 605p 0        800p 0 803p cval 805p 0        1000p 0 1003p 0 1005p 0        1200p 0 1203p 0 1205p 0        1400p 0 1403p cval 1405p 0)
* * I_s0 0 I_s0 pwl(0 0 170p 0 173p cval 175p 0     270p 0 273p cval 275p 0      370p 0 373p 0 375p 0        470p 0 473p cval 475p 0        570p 0 573p 0 575p 0            670p 0 673p 0 675p 0            770p 0 773p cval 775p 0)
* I_z0 0 I_z0 pwl(0 0 200p 0 203p 0 205p 0       400p 0 403p 0 405p 0        600p 0 603p cval 605p 0        800p 0 803p 0 805p 0        1000p 0 1003p cval 1005p 0        1200p 0 1203p cval 1205p 0        1400p 0 1403p cval 1405p 0)


*S = 0 - Select A
*S = 1 - Select B


*A 0
*B   1
*Cin 1

*Expected:
*S 0
*Co 1

* A   0 0 0 1 1 1 1
* B   0 1 1 0 0 1 1
* Ci  1 0 1 0 1 0 1
* S   1 1 0 1 0 0 1
* Cot 0 0 1 0 1 1 1


.tran 0.25p 1600p 0 0.05p

Xsrc_a0 LSmitll_DCSFQ i_a0 src_a0
Xsrc_b0 LSmitll_DCSFQ i_b0 src_b0
Xsrc_ci LSmitll_DCSFQ i_ci src_ci
Xsrc_s0 LSmitll_DCSFQ i_s0 src_s0
Xsrc_z0 LSmitll_DCSFQ i_z0 src_z0

Xload_a0 LSMITLL_JTL src_a0 A0
Xload_b0 LSMITLL_JTL src_b0 B0
Xload_c0 LSMITLL_JTL src_ci Cin
Xload_s0 LSMITLL_JTL src_s0 S_BASE
Xload_z0 LSMITLL_JTL src_z0 Carry_BASE

*For Reference to confirm it is working correctly.
R_QS S_BASE 0 4
R_Cout Carry_BASE 0 4


XDUT DSFQ_ADDDER A0 B0 Cin Sout Cout

* .print p(S_BASE) p(Carry_BASE) p(Sout)  p(CarryOut) p(R3.xdut) p(C3.xdut)
.print p(Sout) p(A0) p(B0) p(Cin) p(Cout)

* .print p(Sout)  p(CarryOut) p(R3.xdut) p(C3.xdut) p(R5.xdut) p(C4.xdut) p(A3.xor1.xdut) p(B3.xor1.xdut)
*  .print p(S_BASE) p(Carry_BASE) p(S)  p(Cout) p(AND1) p(XOR1b) p(AND2) p(C2) p(XOR1b) p(C1)

XCOUT LSMITLL_JTL Cout Carryout
R_Carry Carryout 0 2
XLOAD LSMITLL_JTL S Sout
R_out Sout 0 2

.end