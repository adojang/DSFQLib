.subckt DSFQ_MUX D0 D1 S QQ

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)

.param B2 = 0.8
.param Q2 = 0.8
* .param A2 = 0.8
.param A2 = 0.78
* .param A1 = 3.35
.param A1 = 2
B_x2   B2   	0   	 jjmit area=B2
B_xQ2  	Q2x   	0   	 jjmit area=Q2
B_xA2  	A2   	0   	 jjmit area=A2
B_xA1   A1   	0   	 jjmit area=A1

* XSPLITA LSMITLL_SPLIT1 D0 A1x CLKx
* XSPLITB LSMITLL_SPLITm D1 B1x B1x
* XSPLITS LSMITLL_SPLITm S S1x B2x

* XCJTLA1 LSMITLL_JTLm A1x A1
* XCJTLA2 LSMITLL_JTLm A2x A2
* XCJTLCLK LSMITLL_JTLm CLKx CLK
* XCJTLS1 LSMITLL_JTLm S1x S1
* XCJTLB1 LSMITLL_JTLm B1x B1
* XCJTLB2 LSMITLL_JTLm B2x B2

* XQ1 LSMITLL_JTLm Q1x Q1
* XQ2 LSMITLL_JTLm Q2x Q2


* XAND1   DSFQ_ANDm   A1 A2 Q1x
* XAND2   DSFQ_ANDm   B1 B2 Q2x
* XNOT    DSFQ_NOT S1 CLK CLK A2x
* XOR     DSFQ_ORm    Q1 Q2 QQ



*********************** OR GATE ************************
*OR

LC_OR1_1 Q1 a_OR1 0
LC_OR1_2 Q2 b_OR1 0
LC_OR1_3 QQ Q_OR1 0

* .subckt DSFQ_OR1 a_OR1 b_OR1 q_OR1
.model jjmit_OR1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
*Confluence Buffer A
.param l1_OR1 = 2e-12
.param b1_OR1 = 1.37211310e+00
.param b3_OR1 = 2.77209629e+00
.param b4_OR1 = 3.78734058e-01

* AND GATE LOOP
.param l4_OR1 = 1.22182342e-12
.param b7_OR1 = 1.19265113e+00
.param b9_OR1 = 5.40924075e-01
.param l7_OR1 = 1.62539785e-13
.param r1_OR1 = 1.09745275e+01
.param r2_OR1 = 5.58089917e-01
.param l5_OR1 = 5.61756493e-13

* Output Stage
.param b8_OR1 = 7.09413113e-01
.param i1_OR1 = 3.23631555e-04
.param l3_OR1 = 2e-12
.param l6_OR1 = 3.06315548e-12

*Confluence Buffer B
.param l2_OR1 = L1_OR1
.param b2_OR1 = B1_OR1
.param b5_OR1 = B3_OR1
.param b6_OR1 = B4_OR1

*Parasitics
.param lp1_OR1 = 0.2e-12
.param lp2_OR1 = 0.2e-12
.param lp3_OR1 = 0.2e-12
.param lp4_OR1 = 0.2e-12

* Back Annotated .cir file from KiCad
b1_OR1 3_OR1 1_OR1 jjmit_OR1 area=b1_OR1
b2_OR1 4_OR1 2_OR1 jjmit_OR1 area=b2_OR1
b3_OR1 3_OR1 10_OR1 jjmit_OR1 area=b3_OR1
b4_OR1 5_OR1 3_OR1 jjmit_OR1 area=b4_OR1
b5_OR1 4_OR1 10_OR1 jjmit_OR1 area=b5_OR1
b6_OR1 6_OR1 4_OR1 jjmit_OR1 area=b6_OR1
b7_OR1 24_OR1 20_OR1 jjmit_OR1 area=b7_OR1
b8_OR1 30_OR1 31_OR1 jjmit_OR1 area=b8_OR1
b9_OR1 24_OR1 23_OR1 jjmit_OR1 area=b9_OR1
i1_OR1 0 10_OR1 pwl(0 0 5p i1_OR1)
l1_OR1 a_OR1 1_OR1 l1_OR1
l2_OR1 b_OR1 2_OR1 l2_OR1
l3_OR1 10_OR1 30_OR1 l3_OR1
l4_OR1 30_OR1 20_OR1 l4_OR1
l5_OR1 21_OR1 24_OR1 l5_OR1
l6_OR1 30_OR1 q_OR1 l6_OR1
l7_OR1 22_OR1 23_OR1 l7_OR1
lp1_OR1 5_OR1 0 lp1_OR1
lp2_OR1 6_OR1 0 lp2_OR1
lp3_OR1 24_OR1 0 lp3_OR1
lp4_OR1 31_OR1 0 lp4_OR1
r1_OR1 21_OR1 20_OR1 r1_OR1
r2_OR1 22_OR1 20_OR1 r2_OR1



******************************** AND CELLS ************************************

*AND1
LC_and1_1 A1 a_and1 0
LC_and1_2 A2 b_and1 0
LC_and1_3 Q1x Q_and1 0

.param b1_and1 = 1.39878486e+00
.param bd1_and1 = 1.38855937e+00
.param l1_and1 = 1.64204687e-12
.param rd1_and1 = 6.00718616e-01
.param i1_and1 = 1.54457273e-05
.param b3_and1 = 1.51517089e+00
.param l3_and1 = 2e-12
.param rh1_and1 = 4.76237371e+00
.param ldp1_and1 = 1e-12
.param b2_and1 = b1_and1
.param bd2_and1 = bd1_and1
.param l2_and1 = l1_and1
.param ldp2_and1 = ldp1_and1
.param rd2_and1 = rd1_and1
.param lp1_and1 = 0.2e-12
.param lhp1_and1 = 1e-12
.param lhp2_and1 = lhp1_and1
.param rh2_and1 = rh1_and1

.model jjmit_and1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

b1_and1 30_and1 10_and1 jjmit_and1 area=b1_and1
b2_and1 30_and1 20_and1 jjmit_and1 area=b2_and1
b3_and1 31_and1 30_and1 jjmit_and1 area=b3_and1
bd1_and1 30_and1 12_and1 jjmit_and1 area=bd1_and1
bd2_and1 30_and1 22_and1 jjmit_and1 area=bd2_and1
i1_and1 0 30_and1 pwl(0 0 5p i1_and1)
l1_and1 A_and1 10_and1 l1_and1
l2_and1 B_and1 20_and1 l2_and1
l3_and1 30_and1 Q_and1 l3_and1
ldp1_and1 11_and1 12_and1 ldp1_and1
ldp2_and1 21_and1 22_and1 ldp2_and1
lhp1_and1 13_and1 30_and1 lhp1_and1
lhp2_and1 23_and1 30_and1 lhp2_and1
lp1_and1 31_and1 0 lp1_and1
rd1_and1 11_and1 10_and1 rd1_and1
rd2_and1 21_and1 20_and1 rd2_and1
rh1_and1 13_and1 10_and1 rh1_and1
rh2_and1 23_and1 20_and1 rh2_and1

*AND2
LC_AND2_1 B1 a_AND2 0
LC_AND2_2 B2 b_AND2 0
LC_AND2_3 Q2x Q_AND2 0

.param b1_AND2 = 1.39878486e+00
.param bd1_AND2 = 1.38855937e+00
.param l1_AND2 = 1.64204687e-12
.param rd1_AND2 = 6.00718616e-01
.param i1_AND2 = 1.54457273e-05
.param b3_AND2 = 1.51517089e+00
.param l3_AND2 = 2e-12
.param rh1_AND2 = 4.76237371e+00
.param ldp1_AND2 = 1e-12
.param b2_AND2 = b1_AND2
.param bd2_AND2 = bd1_AND2
.param l2_AND2 = l1_AND2
.param ldp2_AND2 = ldp1_AND2
.param rd2_AND2 = rd1_AND2
.param lp1_AND2 = 0.2e-12
.param lhp1_AND2 = 1e-12
.param lhp2_AND2 = lhp1_AND2
.param rh2_AND2 = rh1_AND2

.model jjmit_AND2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

b1_AND2 30_AND2 10_AND2 jjmit_AND2 area=b1_AND2
b2_AND2 30_AND2 20_AND2 jjmit_AND2 area=b2_AND2
b3_AND2 31_AND2 30_AND2 jjmit_AND2 area=b3_AND2
bd1_AND2 30_AND2 12_AND2 jjmit_AND2 area=bd1_AND2
bd2_AND2 30_AND2 22_AND2 jjmit_AND2 area=bd2_AND2
i1_AND2 0 30_AND2 pwl(0 0 5p i1_AND2)
l1_AND2 A_AND2 10_AND2 l1_AND2
l2_AND2 B_AND2 20_AND2 l2_AND2
l3_AND2 30_AND2 Q_AND2 l3_AND2
ldp1_AND2 11_AND2 12_AND2 ldp1_AND2
ldp2_AND2 21_AND2 22_AND2 ldp2_AND2
lhp1_AND2 13_AND2 30_AND2 lhp1_AND2
lhp2_AND2 23_AND2 30_AND2 lhp2_AND2
lp1_AND2 31_AND2 0 lp1_AND2
rd1_AND2 11_AND2 10_AND2 rd1_AND2
rd2_AND2 21_AND2 20_AND2 rd2_AND2
rh1_AND2 13_AND2 10_AND2 rh1_AND2
rh2_AND2 23_AND2 20_AND2 rh2_AND2






*****JTL CELLS ***********************************************
*JTLA1
LC_JTLA1_1 A1x a_JTLA1 0
LC_JTLA1_2 A1 q_JTLA1 0

.model jjmit_JTLA1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLA1 = 2.0678e-15
.param B0_JTLA1 = 1
.param Ic0_JTLA1 = 1.0000e-04
.param IcRs_JTLA1 = 6.8599e-04
.param B0Rs_JTLA1 = 6.8599
.param Rsheet_JTLA1 = 2
.param Lsheet_JTLA1 = 1.1300e-12
.param LP_JTLA1 = 2.0000e-13
.param IC_JTLA1 = 2.5000
.param Lptl_JTLA1 = 2.0000e-12
.param LB_JTLA1 = 2.0000e-12
.param BiasCoef_JTLA1 = 0.7000
.param B1_JTLA1 = 2.5000
.param B2_JTLA1 = 2.5000
.param IB1_JTLA1 = 3.5000e-04
.param LB1_JTLA1 = 2.0000e-12
.param L1_JTLA1 = 2.0678e-12
.param L2_JTLA1 = 2.0678e-12
.param L3_JTLA1 = 2.0678e-12
.param L4_JTLA1 = 2.0678e-12
.param RB1_JTLA1 = 2.7440
.param RB2_JTLA1 = 2.7440
.param LRB1_JTLA1 = 1.7503e-12
.param LRB2_JTLA1 = 1.7503e-12
.param LP1_JTLA1 = 2.0000e-13
.param LP2_JTLA1 = 2.0000e-13

B1_JTLA1 1_JTLA1 2_JTLA1 jjmit_JTLA1 area=B1_JTLA1
B2_JTLA1 6_JTLA1 7_JTLA1 jjmit_JTLA1 area=B2_JTLA1
IB1_JTLA1 0 5_JTLA1 pwl(0 0 5p IB1_JTLA1)
L1_JTLA1 a_JTLA1 1_JTLA1 2.082E-12
L2_JTLA1 1_JTLA1 4_JTLA1 2.06E-12
L3_JTLA1 4_JTLA1 6_JTLA1 2.067E-12
L4_JTLA1 6_JTLA1 q_JTLA1 2.075E-12
LP1_JTLA1 2_JTLA1 0 4.998E-13
LP2_JTLA1 7_JTLA1 0 5.011E-13
LB1_JTLA1 5_JTLA1 4_JTLA1 LB1_JTLA1
RB1_JTLA1 1_JTLA1 3_JTLA1 RB1_JTLA1
RB2_JTLA1 6_JTLA1 8_JTLA1 RB2_JTLA1
LRB1_JTLA1 3_JTLA1 0 LRB1_JTLA1
LRB2_JTLA1 8_JTLA1 0 LRB2_JTLA1

*JTLA2
LC_JTLA2_1 A2x a_JTLA2 0
LC_JTLA2_2 A2 q_JTLA2 0

.model jjmit_JTLA2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLA2 = 2.0678e-15
.param B0_JTLA2 = 1
.param Ic0_JTLA2 = 1.0000e-04
.param IcRs_JTLA2 = 6.8599e-04
.param B0Rs_JTLA2 = 6.8599
.param Rsheet_JTLA2 = 2
.param Lsheet_JTLA2 = 1.1300e-12
.param LP_JTLA2 = 2.0000e-13
.param IC_JTLA2 = 2.5000
.param Lptl_JTLA2 = 2.0000e-12
.param LB_JTLA2 = 2.0000e-12
.param BiasCoef_JTLA2 = 0.7000
.param B1_JTLA2 = 2.5000
.param B2_JTLA2 = 2.5000
.param IB1_JTLA2 = 3.5000e-04
.param LB1_JTLA2 = 2.0000e-12
.param L1_JTLA2 = 2.0678e-12
.param L2_JTLA2 = 2.0678e-12
.param L3_JTLA2 = 2.0678e-12
.param L4_JTLA2 = 2.0678e-12
.param RB1_JTLA2 = 2.7440
.param RB2_JTLA2 = 2.7440
.param LRB1_JTLA2 = 1.7503e-12
.param LRB2_JTLA2 = 1.7503e-12
.param LP1_JTLA2 = 2.0000e-13
.param LP2_JTLA2 = 2.0000e-13

B1_JTLA2 1_JTLA2 2_JTLA2 jjmit_JTLA2 area=B1_JTLA2
B2_JTLA2 6_JTLA2 7_JTLA2 jjmit_JTLA2 area=B2_JTLA2
IB1_JTLA2 0 5_JTLA2 pwl(0 0 5p IB1_JTLA2)
L1_JTLA2 a_JTLA2 1_JTLA2 2.082E-12
L2_JTLA2 1_JTLA2 4_JTLA2 2.06E-12
L3_JTLA2 4_JTLA2 6_JTLA2 2.067E-12
L4_JTLA2 6_JTLA2 q_JTLA2 2.075E-12
LP1_JTLA2 2_JTLA2 0 4.998E-13
LP2_JTLA2 7_JTLA2 0 5.011E-13
LB1_JTLA2 5_JTLA2 4_JTLA2 LB1_JTLA2
RB1_JTLA2 1_JTLA2 3_JTLA2 RB1_JTLA2
RB2_JTLA2 6_JTLA2 8_JTLA2 RB2_JTLA2
LRB1_JTLA2 3_JTLA2 0 LRB1_JTLA2
LRB2_JTLA2 8_JTLA2 0 LRB2_JTLA2

*JTLCLK
LC_JTLCLK_1 CLKx a_JTLCLK 0
LC_JTLCLK_2 CLK q_JTLCLK 0

.model jjmit_JTLCLK jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLCLK = 2.0678e-15
.param B0_JTLCLK = 1
.param Ic0_JTLCLK = 1.0000e-04
.param IcRs_JTLCLK = 6.8599e-04
.param B0Rs_JTLCLK = 6.8599
.param Rsheet_JTLCLK = 2
.param Lsheet_JTLCLK = 1.1300e-12
.param LP_JTLCLK = 2.0000e-13
.param IC_JTLCLK = 2.5000
.param Lptl_JTLCLK = 2.0000e-12
.param LB_JTLCLK = 2.0000e-12
.param BiasCoef_JTLCLK = 0.7000
.param B1_JTLCLK = 2.5000
.param B2_JTLCLK = 2.5000
.param IB1_JTLCLK = 3.5000e-04
.param LB1_JTLCLK = 2.0000e-12
.param L1_JTLCLK = 2.0678e-12
.param L2_JTLCLK = 2.0678e-12
.param L3_JTLCLK = 2.0678e-12
.param L4_JTLCLK = 2.0678e-12
.param RB1_JTLCLK = 2.7440
.param RB2_JTLCLK = 2.7440
.param LRB1_JTLCLK = 1.7503e-12
.param LRB2_JTLCLK = 1.7503e-12
.param LP1_JTLCLK = 2.0000e-13
.param LP2_JTLCLK = 2.0000e-13

B1_JTLCLK 1_JTLCLK 2_JTLCLK jjmit_JTLCLK area=B1_JTLCLK
B2_JTLCLK 6_JTLCLK 7_JTLCLK jjmit_JTLCLK area=B2_JTLCLK
IB1_JTLCLK 0 5_JTLCLK pwl(0 0 5p IB1_JTLCLK)
L1_JTLCLK a_JTLCLK 1_JTLCLK 2.082E-12
L2_JTLCLK 1_JTLCLK 4_JTLCLK 2.06E-12
L3_JTLCLK 4_JTLCLK 6_JTLCLK 2.067E-12
L4_JTLCLK 6_JTLCLK q_JTLCLK 2.075E-12
LP1_JTLCLK 2_JTLCLK 0 4.998E-13
LP2_JTLCLK 7_JTLCLK 0 5.011E-13
LB1_JTLCLK 5_JTLCLK 4_JTLCLK LB1_JTLCLK
RB1_JTLCLK 1_JTLCLK 3_JTLCLK RB1_JTLCLK
RB2_JTLCLK 6_JTLCLK 8_JTLCLK RB2_JTLCLK
LRB1_JTLCLK 3_JTLCLK 0 LRB1_JTLCLK
LRB2_JTLCLK 8_JTLCLK 0 LRB2_JTLCLK


*JTLS1
LC_JTLS1_1 S1x a_JTLS1 0
LC_JTLS1_2 S1 q_JTLS1 0

.model jjmit_JTLS1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLS1 = 2.0678e-15
.param B0_JTLS1 = 1
.param Ic0_JTLS1 = 1.0000e-04
.param IcRs_JTLS1 = 6.8599e-04
.param B0Rs_JTLS1 = 6.8599
.param Rsheet_JTLS1 = 2
.param Lsheet_JTLS1 = 1.1300e-12
.param LP_JTLS1 = 2.0000e-13
.param IC_JTLS1 = 2.5000
.param Lptl_JTLS1 = 2.0000e-12
.param LB_JTLS1 = 2.0000e-12
.param BiasCoef_JTLS1 = 0.7000
.param B1_JTLS1 = 2.5000
.param B2_JTLS1 = 2.5000
.param IB1_JTLS1 = 3.5000e-04
.param LB1_JTLS1 = 2.0000e-12
.param L1_JTLS1 = 2.0678e-12
.param L2_JTLS1 = 2.0678e-12
.param L3_JTLS1 = 2.0678e-12
.param L4_JTLS1 = 2.0678e-12
.param RB1_JTLS1 = 2.7440
.param RB2_JTLS1 = 2.7440
.param LRB1_JTLS1 = 1.7503e-12
.param LRB2_JTLS1 = 1.7503e-12
.param LP1_JTLS1 = 2.0000e-13
.param LP2_JTLS1 = 2.0000e-13

B1_JTLS1 1_JTLS1 2_JTLS1 jjmit_JTLS1 area=B1_JTLS1
B2_JTLS1 6_JTLS1 7_JTLS1 jjmit_JTLS1 area=B2_JTLS1
IB1_JTLS1 0 5_JTLS1 pwl(0 0 5p IB1_JTLS1)
L1_JTLS1 a_JTLS1 1_JTLS1 2.082E-12
L2_JTLS1 1_JTLS1 4_JTLS1 2.06E-12
L3_JTLS1 4_JTLS1 6_JTLS1 2.067E-12
L4_JTLS1 6_JTLS1 q_JTLS1 2.075E-12
LP1_JTLS1 2_JTLS1 0 4.998E-13
LP2_JTLS1 7_JTLS1 0 5.011E-13
LB1_JTLS1 5_JTLS1 4_JTLS1 LB1_JTLS1
RB1_JTLS1 1_JTLS1 3_JTLS1 RB1_JTLS1
RB2_JTLS1 6_JTLS1 8_JTLS1 RB2_JTLS1
LRB1_JTLS1 3_JTLS1 0 LRB1_JTLS1
LRB2_JTLS1 8_JTLS1 0 LRB2_JTLS1

*JTLB1
LC_JTLB1_1 B1x a_JTLB1 0
LC_JTLB1_2 B1 q_JTLB1 0

.model jjmit_JTLB1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLB1 = 2.0678e-15
.param B0_JTLB1 = 1
.param Ic0_JTLB1 = 1.0000e-04
.param IcRs_JTLB1 = 6.8599e-04
.param B0Rs_JTLB1 = 6.8599
.param Rsheet_JTLB1 = 2
.param Lsheet_JTLB1 = 1.1300e-12
.param LP_JTLB1 = 2.0000e-13
.param IC_JTLB1 = 2.5000
.param Lptl_JTLB1 = 2.0000e-12
.param LB_JTLB1 = 2.0000e-12
.param BiasCoef_JTLB1 = 0.7000
.param B1_JTLB1 = 2.5000
.param B2_JTLB1 = 2.5000
.param IB1_JTLB1 = 3.5000e-04
.param LB1_JTLB1 = 2.0000e-12
.param L1_JTLB1 = 2.0678e-12
.param L2_JTLB1 = 2.0678e-12
.param L3_JTLB1 = 2.0678e-12
.param L4_JTLB1 = 2.0678e-12
.param RB1_JTLB1 = 2.7440
.param RB2_JTLB1 = 2.7440
.param LRB1_JTLB1 = 1.7503e-12
.param LRB2_JTLB1 = 1.7503e-12
.param LP1_JTLB1 = 2.0000e-13
.param LP2_JTLB1 = 2.0000e-13

B1_JTLB1 1_JTLB1 2_JTLB1 jjmit_JTLB1 area=B1_JTLB1
B2_JTLB1 6_JTLB1 7_JTLB1 jjmit_JTLB1 area=B2_JTLB1
IB1_JTLB1 0 5_JTLB1 pwl(0 0 5p IB1_JTLB1)
L1_JTLB1 a_JTLB1 1_JTLB1 2.082E-12
L2_JTLB1 1_JTLB1 4_JTLB1 2.06E-12
L3_JTLB1 4_JTLB1 6_JTLB1 2.067E-12
L4_JTLB1 6_JTLB1 q_JTLB1 2.075E-12
LP1_JTLB1 2_JTLB1 0 4.998E-13
LP2_JTLB1 7_JTLB1 0 5.011E-13
LB1_JTLB1 5_JTLB1 4_JTLB1 LB1_JTLB1
RB1_JTLB1 1_JTLB1 3_JTLB1 RB1_JTLB1
RB2_JTLB1 6_JTLB1 8_JTLB1 RB2_JTLB1
LRB1_JTLB1 3_JTLB1 0 LRB1_JTLB1
LRB2_JTLB1 8_JTLB1 0 LRB2_JTLB1

*JTLB2
LC_JTLB2_1 B2x a_JTLB2 0
LC_JTLB2_2 B2 q_JTLB2 0

.model jjmit_JTLB2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLB2 = 2.0678e-15
.param B0_JTLB2 = 1
.param Ic0_JTLB2 = 1.0000e-04
.param IcRs_JTLB2 = 6.8599e-04
.param B0Rs_JTLB2 = 6.8599
.param Rsheet_JTLB2 = 2
.param Lsheet_JTLB2 = 1.1300e-12
.param LP_JTLB2 = 2.0000e-13
.param IC_JTLB2 = 2.5000
.param Lptl_JTLB2 = 2.0000e-12
.param LB_JTLB2 = 2.0000e-12
.param BiasCoef_JTLB2 = 0.7000
.param B1_JTLB2 = 2.5000
.param B2_JTLB2 = 2.5000
.param IB1_JTLB2 = 3.5000e-04
.param LB1_JTLB2 = 2.0000e-12
.param L1_JTLB2 = 2.0678e-12
.param L2_JTLB2 = 2.0678e-12
.param L3_JTLB2 = 2.0678e-12
.param L4_JTLB2 = 2.0678e-12
.param RB1_JTLB2 = 2.7440
.param RB2_JTLB2 = 2.7440
.param LRB1_JTLB2 = 1.7503e-12
.param LRB2_JTLB2 = 1.7503e-12
.param LP1_JTLB2 = 2.0000e-13
.param LP2_JTLB2 = 2.0000e-13

B1_JTLB2 1_JTLB2 2_JTLB2 jjmit_JTLB2 area=B1_JTLB2
B2_JTLB2 6_JTLB2 7_JTLB2 jjmit_JTLB2 area=B2_JTLB2
IB1_JTLB2 0 5_JTLB2 pwl(0 0 5p IB1_JTLB2)
L1_JTLB2 a_JTLB2 1_JTLB2 2.082E-12
L2_JTLB2 1_JTLB2 4_JTLB2 2.06E-12
L3_JTLB2 4_JTLB2 6_JTLB2 2.067E-12
L4_JTLB2 6_JTLB2 q_JTLB2 2.075E-12
LP1_JTLB2 2_JTLB2 0 4.998E-13
LP2_JTLB2 7_JTLB2 0 5.011E-13
LB1_JTLB2 5_JTLB2 4_JTLB2 LB1_JTLB2
RB1_JTLB2 1_JTLB2 3_JTLB2 RB1_JTLB2
RB2_JTLB2 6_JTLB2 8_JTLB2 RB2_JTLB2
LRB1_JTLB2 3_JTLB2 0 LRB1_JTLB2
LRB2_JTLB2 8_JTLB2 0 LRB2_JTLB2


*JTLQ1
LC_JTLQ1_1 Q1x a_JTLQ1 0
LC_JTLQ1_2 Q1 q_JTLQ1 0

.model jjmit_JTLQ1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLQ1 = 2.0678e-15
.param B0_JTLQ1 = 1
.param Ic0_JTLQ1 = 1.0000e-04
.param IcRs_JTLQ1 = 6.8599e-04
.param B0Rs_JTLQ1 = 6.8599
.param Rsheet_JTLQ1 = 2
.param Lsheet_JTLQ1 = 1.1300e-12
.param LP_JTLQ1 = 2.0000e-13
.param IC_JTLQ1 = 2.5000
.param Lptl_JTLQ1 = 2.0000e-12
.param LB_JTLQ1 = 2.0000e-12
.param BiasCoef_JTLQ1 = 0.7000
.param B1_JTLQ1 = 2.5000
.param B2_JTLQ1 = 2.5000
.param IB1_JTLQ1 = 3.5000e-04
.param LB1_JTLQ1 = 2.0000e-12
.param L1_JTLQ1 = 2.0678e-12
.param L2_JTLQ1 = 2.0678e-12
.param L3_JTLQ1 = 2.0678e-12
.param L4_JTLQ1 = 2.0678e-12
.param RB1_JTLQ1 = 2.7440
.param RB2_JTLQ1 = 2.7440
.param LRB1_JTLQ1 = 1.7503e-12
.param LRB2_JTLQ1 = 1.7503e-12
.param LP1_JTLQ1 = 2.0000e-13
.param LP2_JTLQ1 = 2.0000e-13

B1_JTLQ1 1_JTLQ1 2_JTLQ1 jjmit_JTLQ1 area=B1_JTLQ1
B2_JTLQ1 6_JTLQ1 7_JTLQ1 jjmit_JTLQ1 area=B2_JTLQ1
IB1_JTLQ1 0 5_JTLQ1 pwl(0 0 5p IB1_JTLQ1)
L1_JTLQ1 a_JTLQ1 1_JTLQ1 2.082E-12
L2_JTLQ1 1_JTLQ1 4_JTLQ1 2.06E-12
L3_JTLQ1 4_JTLQ1 6_JTLQ1 2.067E-12
L4_JTLQ1 6_JTLQ1 q_JTLQ1 2.075E-12
LP1_JTLQ1 2_JTLQ1 0 4.998E-13
LP2_JTLQ1 7_JTLQ1 0 5.011E-13
LB1_JTLQ1 5_JTLQ1 4_JTLQ1 LB1_JTLQ1
RB1_JTLQ1 1_JTLQ1 3_JTLQ1 RB1_JTLQ1
RB2_JTLQ1 6_JTLQ1 8_JTLQ1 RB2_JTLQ1
LRB1_JTLQ1 3_JTLQ1 0 LRB1_JTLQ1
LRB2_JTLQ1 8_JTLQ1 0 LRB2_JTLQ1

*JTLQ2
LC_JTLQ2_1 Q2x a_JTLQ2 0
LC_JTLQ2_2 Q2 q_JTLQ2 0

.model jjmit_JTLQ2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLQ2 = 2.0678e-15
.param B0_JTLQ2 = 1
.param Ic0_JTLQ2 = 1.0000e-04
.param IcRs_JTLQ2 = 6.8599e-04
.param B0Rs_JTLQ2 = 6.8599
.param Rsheet_JTLQ2 = 2
.param Lsheet_JTLQ2 = 1.1300e-12
.param LP_JTLQ2 = 2.0000e-13
.param IC_JTLQ2 = 2.5000
.param Lptl_JTLQ2 = 2.0000e-12
.param LB_JTLQ2 = 2.0000e-12
.param BiasCoef_JTLQ2 = 0.7000
.param B1_JTLQ2 = 2.5000
.param B2_JTLQ2 = 2.5000
.param IB1_JTLQ2 = 3.5000e-04
.param LB1_JTLQ2 = 2.0000e-12
.param L1_JTLQ2 = 2.0678e-12
.param L2_JTLQ2 = 2.0678e-12
.param L3_JTLQ2 = 2.0678e-12
.param L4_JTLQ2 = 2.0678e-12
.param RB1_JTLQ2 = 2.7440
.param RB2_JTLQ2 = 2.7440
.param LRB1_JTLQ2 = 1.7503e-12
.param LRB2_JTLQ2 = 1.7503e-12
.param LP1_JTLQ2 = 2.0000e-13
.param LP2_JTLQ2 = 2.0000e-13

B1_JTLQ2 1_JTLQ2 2_JTLQ2 jjmit_JTLQ2 area=B1_JTLQ2
B2_JTLQ2 6_JTLQ2 7_JTLQ2 jjmit_JTLQ2 area=B2_JTLQ2
IB1_JTLQ2 0 5_JTLQ2 pwl(0 0 5p IB1_JTLQ2)
L1_JTLQ2 a_JTLQ2 1_JTLQ2 2.082E-12
L2_JTLQ2 1_JTLQ2 4_JTLQ2 2.06E-12
L3_JTLQ2 4_JTLQ2 6_JTLQ2 2.067E-12
L4_JTLQ2 6_JTLQ2 q_JTLQ2 2.075E-12
LP1_JTLQ2 2_JTLQ2 0 4.998E-13
LP2_JTLQ2 7_JTLQ2 0 5.011E-13
LB1_JTLQ2 5_JTLQ2 4_JTLQ2 LB1_JTLQ2
RB1_JTLQ2 1_JTLQ2 3_JTLQ2 RB1_JTLQ2
RB2_JTLQ2 6_JTLQ2 8_JTLQ2 RB2_JTLQ2
LRB1_JTLQ2 3_JTLQ2 0 LRB1_JTLQ2
LRB2_JTLQ2 8_JTLQ2 0 LRB2_JTLQ2




*** SPLIT CELLS********************************************************************************************************************************

LC_split1_1 D0 a_split1 0
LC_split1_2 A1x q0_split1 0
LC_split1_3 CLKx q1_split1 0
.model jjmit_split1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_split1 = 2.0678e-15
.param B0_split1 = 1
.param Ic0_split1 = 1.0000e-04
.param IcRs_split1 = 6.8599e-04
.param B0Rs_split1 = 6.8599
.param Rsheet_split1 = 2
.param Lsheet_split1 = 1.1300e-12
.param LP_split1 = 2.0000e-13
.param IC_split1 = 2.5000
.param Lptl_split1 = 2.0000e-12
.param LB_split1 = 2.0000e-12
.param BiasCoef_split1 = 0.7000
.param RD_split1 = 1.3600
.param B1_split1 = 2.5000
.param B2_split1 = 3
.param B3_split1 = 2.5000
.param B4_split1 = 2.5000
.param IB1_split1 = 1.7500e-04
.param IB2_split1 = 2.8000e-04
.param IB3_split1 = 1.7500e-04
.param IB4_split1 = 1.7500e-04
.param L1_split1 = 2.0000e-12
.param L2_split1 = 4.1357e-12
.param L3_split1 = 1.7232e-12
.param L4_split1 = 1.7232e-12
.param L5_split1 = 2.0000e-12
.param L6_split1 = 1.7232e-12
.param L7_split1 = 2.0000e-12
.param RB1_split1 = 2.7440
.param RB2_split1 = 2.2866
.param RB3_split1 = 2.7440
.param RB4_split1 = 2.7440
.param LRB1_split1 = 1.5503e-12
.param LRB2_split1 = 1.2919e-12
.param LRB3_split1 = 1.5503e-12
.param LRB4_split1 = 1.5503e-12

IB1_split1 0 3_split1 pwl(0 0 5p IB1_split1)
IB2_split1 0 6_split1 pwl(0 0 5p IB2_split1)
IB3_split1 0 10_split1 pwl(0 0 5p IB3_split1)
IB4_split1 0 13_split1 pwl(0 0 5p IB4_split1)
LB1_split1 3_split1 1_split1 9.175E-13
LB2_split1 6_split1 4_split1 7.666E-13
LB3_split1 10_split1 8_split1 1.928E-12
LB4_split1 13_split1 11_split1 8.786E-13

B1_split1 1_split1 2_split1 jjmit_split1 area=B1_split1
B2_split1 4_split1 5_split1 jjmit_split1 area=B2_split1
B3_split1 8_split1 9_split1 jjmit_split1 area=B3_split1
B4_split1 11_split1 12_split1 jjmit_split1 area=B4_split1
L1_split1 a_split1 1_split1 2.063E-12
L2_split1 1_split1 4_split1 3.637E-12
L3_split1 4_split1 7_split1 1.278E-12
L4_split1 7_split1 8_split1 1.305E-12
L5_split1 8_split1 q0_split1 2.05E-12
L6_split1 7_split1 11_split1 1.315E-12
L7_split1 11_split1 q1_split1 2.06E-12

LP1_split1 2_split1 0 4.676E-13
LP2_split1 5_split1 0 4.498E-13
LP3_split1 9_split1 0 5.183E-13
LP4_split1 12_split1 0 4.639E-13
RB1_split1 1_split1 101_split1 RB1_split1
LRB1_split1 101_split1 0 LRB1_split1
RB2_split1 4_split1 104_split1 RB2_split1
LRB2_split1 104_split1 0 LRB2_split1
RB3_split1 8_split1 108_split1 RB3_split1
LRB3_split1 108_split1 0 LRB3_split1
RB4_split1 11_split1 111_split1 RB4_split1
LRB4_split1 111_split1 0 LRB4_split1



*SPLIT2



LC_split2_1 D1 a_split2 0
LC_split2_2 B1x q0_split2 0
LC_split2_3 B1x q1_split2 0
.model jjmit_split2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_split2 = 2.0678e-15
.param B0_split2 = 1
.param Ic0_split2 = 1.0000e-04
.param IcRs_split2 = 6.8599e-04
.param B0Rs_split2 = 6.8599
.param Rsheet_split2 = 2
.param Lsheet_split2 = 1.1300e-12
.param LP_split2 = 2.0000e-13
.param IC_split2 = 2.5000
.param Lptl_split2 = 2.0000e-12
.param LB_split2 = 2.0000e-12
.param BiasCoef_split2 = 0.7000
.param RD_split2 = 1.3600
.param B1_split2 = 2.5000
.param B2_split2 = 3
.param B3_split2 = 2.5000
.param B4_split2 = 2.5000
.param IB1_split2 = 1.7500e-04
.param IB2_split2 = 2.8000e-04
.param IB3_split2 = 1.7500e-04
.param IB4_split2 = 1.7500e-04
.param L1_split2 = 2.0000e-12
.param L2_split2 = 4.1357e-12
.param L3_split2 = 1.7232e-12
.param L4_split2 = 1.7232e-12
.param L5_split2 = 2.0000e-12
.param L6_split2 = 1.7232e-12
.param L7_split2 = 2.0000e-12
.param RB1_split2 = 2.7440
.param RB2_split2 = 2.2866
.param RB3_split2 = 2.7440
.param RB4_split2 = 2.7440
.param LRB1_split2 = 1.5503e-12
.param LRB2_split2 = 1.2919e-12
.param LRB3_split2 = 1.5503e-12
.param LRB4_split2 = 1.5503e-12

IB1_split2 0 3_split2 pwl(0 0 5p IB1_split2)
IB2_split2 0 6_split2 pwl(0 0 5p IB2_split2)
IB3_split2 0 10_split2 pwl(0 0 5p IB3_split2)
IB4_split2 0 13_split2 pwl(0 0 5p IB4_split2)
LB1_split2 3_split2 1_split2 9.175E-13
LB2_split2 6_split2 4_split2 7.666E-13
LB3_split2 10_split2 8_split2 1.928E-12
LB4_split2 13_split2 11_split2 8.786E-13

B1_split2 1_split2 2_split2 jjmit_split2 area=B1_split2
B2_split2 4_split2 5_split2 jjmit_split2 area=B2_split2
B3_split2 8_split2 9_split2 jjmit_split2 area=B3_split2
B4_split2 11_split2 12_split2 jjmit_split2 area=B4_split2
L1_split2 a_split2 1_split2 2.063E-12
L2_split2 1_split2 4_split2 3.637E-12
L3_split2 4_split2 7_split2 1.278E-12
L4_split2 7_split2 8_split2 1.305E-12
L5_split2 8_split2 q0_split2 2.05E-12
L6_split2 7_split2 11_split2 1.315E-12
L7_split2 11_split2 q1_split2 2.06E-12

LP1_split2 2_split2 0 4.676E-13
LP2_split2 5_split2 0 4.498E-13
LP3_split2 9_split2 0 5.183E-13
LP4_split2 12_split2 0 4.639E-13
RB1_split2 1_split2 101_split2 RB1_split2
LRB1_split2 101_split2 0 LRB1_split2
RB2_split2 4_split2 104_split2 RB2_split2
LRB2_split2 104_split2 0 LRB2_split2
RB3_split2 8_split2 108_split2 RB3_split2
LRB3_split2 108_split2 0 LRB3_split2
RB4_split2 11_split2 111_split2 RB4_split2
LRB4_split2 111_split2 0 LRB4_split2

*SPLIT3

LC_split3_1 S a_split3 0
LC_split3_2 S1x q0_split3 0
LC_split3_3 B2x q1_split3 0
.model jjmit_split3 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_split3 = 2.0678e-15
.param B0_split3 = 1
.param Ic0_split3 = 1.0000e-04
.param IcRs_split3 = 6.8599e-04
.param B0Rs_split3 = 6.8599
.param Rsheet_split3 = 2
.param Lsheet_split3 = 1.1300e-12
.param LP_split3 = 2.0000e-13
.param IC_split3 = 2.5000
.param Lptl_split3 = 2.0000e-12
.param LB_split3 = 2.0000e-12
.param BiasCoef_split3 = 0.7000
.param RD_split3 = 1.3600
.param B1_split3 = 2.5000
.param B2_split3 = 3
.param B3_split3 = 2.5000
.param B4_split3 = 2.5000
.param IB1_split3 = 1.7500e-04
.param IB2_split3 = 2.8000e-04
.param IB3_split3 = 1.7500e-04
.param IB4_split3 = 1.7500e-04
.param L1_split3 = 2.0000e-12
.param L2_split3 = 4.1357e-12
.param L3_split3 = 1.7232e-12
.param L4_split3 = 1.7232e-12
.param L5_split3 = 2.0000e-12
.param L6_split3 = 1.7232e-12
.param L7_split3 = 2.0000e-12
.param RB1_split3 = 2.7440
.param RB2_split3 = 2.2866
.param RB3_split3 = 2.7440
.param RB4_split3 = 2.7440
.param LRB1_split3 = 1.5503e-12
.param LRB2_split3 = 1.2919e-12
.param LRB3_split3 = 1.5503e-12
.param LRB4_split3 = 1.5503e-12

IB1_split3 0 3_split3 pwl(0 0 5p IB1_split3)
IB2_split3 0 6_split3 pwl(0 0 5p IB2_split3)
IB3_split3 0 10_split3 pwl(0 0 5p IB3_split3)
IB4_split3 0 13_split3 pwl(0 0 5p IB4_split3)
LB1_split3 3_split3 1_split3 9.175E-13
LB2_split3 6_split3 4_split3 7.666E-13
LB3_split3 10_split3 8_split3 1.928E-12
LB4_split3 13_split3 11_split3 8.786E-13

B1_split3 1_split3 2_split3 jjmit_split3 area=B1_split3
B2_split3 4_split3 5_split3 jjmit_split3 area=B2_split3
B3_split3 8_split3 9_split3 jjmit_split3 area=B3_split3
B4_split3 11_split3 12_split3 jjmit_split3 area=B4_split3
L1_split3 a_split3 1_split3 2.063E-12
L2_split3 1_split3 4_split3 3.637E-12
L3_split3 4_split3 7_split3 1.278E-12
L4_split3 7_split3 8_split3 1.305E-12
L5_split3 8_split3 q0_split3 2.05E-12
L6_split3 7_split3 11_split3 1.315E-12
L7_split3 11_split3 q1_split3 2.06E-12

LP1_split3 2_split3 0 4.676E-13
LP2_split3 5_split3 0 4.498E-13
LP3_split3 9_split3 0 5.183E-13
LP4_split3 12_split3 0 4.639E-13
RB1_split3 1_split3 101_split3 RB1_split3
LRB1_split3 101_split3 0 LRB1_split3
RB2_split3 4_split3 104_split3 RB2_split3
LRB2_split3 104_split3 0 LRB2_split3
RB3_split3 8_split3 108_split3 RB3_split3
LRB3_split3 108_split3 0 LRB3_split3
RB4_split3 11_split3 111_split3 RB4_split3
LRB4_split3 111_split3 0 LRB4_split3


*****************************************************************************************************

*NOT

LC_NOT_1 S1 Ann 0
LC_NOT_2 CLK Bnn 0
LC_NOT_3 CLK Cnn 0
LC_NOT_4 A2x Qnn 0
* .subckt DSFQ_NOT A B C Q
*A is inverting input.
*B and C are inputs for the OR gate.
*Q is output.

* XDSFQ_OR DSFQ_OR B C CLK
* XJTLCLK LSMITLL_JTLi CLK CLK1
* XNOTLS LSMITLL_NOTi A CLK1 Q


LC_NOT_OR_1 Bnn a_NOT_OR 0
LC_NOT_OR_2 Cnn b_NOT_OR 0
LC_NOT_OR_3 CLKnn q_NOT_OR 0
*OR GATE
.model jjmit_NOT_OR jj(rtype=1_NOT_OR, vg=2.8mV_NOT_OR, cap=0.07pF_NOT_OR, r0=160_NOT_OR, rn=16_NOT_OR, icrit=0.1mA_NOT_OR)

*Confluence Buffer A
.param l1_NOT_OR = 0.001e-12
.param b1_NOT_OR = 1.44497758
.param b3_NOT_OR = 5.41067564
.param b4_NOT_OR = 7.95470698

* AND GATE LOOP
.param l4_NOT_OR = 1.22182342e-12
.param b7_NOT_OR = 1.59265113
.param b9_NOT_OR = 5.40924075e-01
.param l7_NOT_OR = 1.62539785e-13
.param r1_NOT_OR = 1.09745275e+01
.param r2_NOT_OR = 5.58089917e-01
.param l5_NOT_OR = 5.61756493e-13

* Output Stage
.param b8_NOT_OR = 4.73543077e-01
.param i1_NOT_OR = 3.40214819e-04
.param l3_NOT_OR = 2e-12
.param l6_NOT_OR = 3.06315548e-12

*Confluence Buffer B
.param l2_NOT_OR = l1_NOT_OR
.param b2_NOT_OR = b1_NOT_OR
.param b5_NOT_OR = b3_NOT_OR
.param b6_NOT_OR = b4_NOT_OR

*Parasitics
.param lp1_NOT_OR = 0.2e-12
.param lp2_NOT_OR = 0.2e-12
.param lp3_NOT_OR = 0.2e-12
.param lp4_NOT_OR = 0.2e-12

* Back Annotated .cir file from KiCad
b1_NOT_OR 3_NOT_OR 1_NOT_OR jjmit_NOT_OR area=b1_NOT_OR
b2_NOT_OR 4_NOT_OR 2_NOT_OR jjmit_NOT_OR area=b2_NOT_OR
b3_NOT_OR 3_NOT_OR 10_NOT_OR jjmit_NOT_OR area=b3_NOT_OR
b4_NOT_OR 5_NOT_OR 3_NOT_OR jjmit_NOT_OR area=b4_NOT_OR
b5_NOT_OR 4_NOT_OR 10_NOT_OR jjmit_NOT_OR area=b5_NOT_OR
b6_NOT_OR 6_NOT_OR 4_NOT_OR jjmit_NOT_OR area=b6_NOT_OR
b7_NOT_OR 24_NOT_OR 20_NOT_OR jjmit_NOT_OR area=b7_NOT_OR
b8_NOT_OR 30_NOT_OR 31_NOT_OR jjmit_NOT_OR area=b8_NOT_OR
b9_NOT_OR 24_NOT_OR 23_NOT_OR jjmit_NOT_OR area=b9_NOT_OR
i1_NOT_OR 0 10_NOT_OR pwl(0 0 5p i1_NOT_OR)
l1_NOT_OR a_NOT_OR 1_NOT_OR l1_NOT_OR
l2_NOT_OR b_NOT_OR 2_NOT_OR l2_NOT_OR
l3_NOT_OR 10_NOT_OR 30_NOT_OR l3_NOT_OR
l4_NOT_OR 30_NOT_OR 20_NOT_OR l4_NOT_OR
l5_NOT_OR 21_NOT_OR 24_NOT_OR l5_NOT_OR
l6_NOT_OR 30_NOT_OR q_NOT_OR l6_NOT_OR
l7_NOT_OR 22_NOT_OR 23_NOT_OR l7_NOT_OR
lp1_NOT_OR 5_NOT_OR 0 lp1_NOT_OR
lp2_NOT_OR 6_NOT_OR 0 lp2_NOT_OR
lp3_NOT_OR 24_NOT_OR 0 lp3_NOT_OR
lp4_NOT_OR 31_NOT_OR 0 lp4_NOT_OR
r1_NOT_OR 21_NOT_OR 20_NOT_OR r1_NOT_OR
r2_NOT_OR 22_NOT_OR 20_NOT_OR r2_NOT_OR

*NOT
LC_NOT_NOT_1 Ann a_NOT1 0
LC_NOT_NOT_2 CLK1nn clk_NOT1 0
LC_NOT_NOT_3 Qnn q_NOT1 0

.model jjmit_NOT1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

.param Phi0_NOT1 = 2.0678e-15
.param B0_NOT1 = 1
.param Ic0_NOT1 = 1.0000e-04
.param IcRs_NOT1 = 6.8599e-04
.param B0Rs_NOT1 = 6.8599
.param Rsheet_NOT1 = 2
.param Lsheet_NOT1 = 1.1300e-12
.param LP_NOT1 = 2.0000e-13
.param IC_NOT1 = 2.5000
.param LB_NOT1 = 2.0000e-12
.param BiasCoef_NOT1 = 0.7000
.param B1_NOT1 = 2.5000
.param B2_NOT1 = 2.5700
.param B3_NOT1 = 1.0700
.param B4_NOT1 = 2.5000
.param B5_NOT1 = 1.3400
.param B6_NOT1 = 3.0300
.param B7_NOT1 = 1.3800
.param B8_NOT1 = 0.8000
.param B9_NOT1 = 2.5000
.param IB1_NOT1 = 1.7500e-04
.param IB2_NOT1 = 8.7000e-05
.param IB3_NOT1 = 2.5700e-04
.param IB4_NOT1 = 1.7500e-04
.param IB5_NOT1 = 1.7500e-04
.param LB1_NOT1 = 2.0000e-12
.param LB2_NOT1 = 2.0000e-12
.param LB3_NOT1 = 2.0000e-12
.param LB4_NOT1 = 2.0000e-12
.param LB5_NOT1 = 2.0000e-12
.param RB1_NOT1 = 2.7440
.param RB2_NOT1 = 2.6692
.param RB3_NOT1 = 6.4111
.param RB4_NOT1 = 2.7440
.param RB5_NOT1 = 5.1193
.param RB6_NOT1 = 2.2640
.param RB7_NOT1 = 4.9709
.param RB8_NOT1 = 8.5749
.param RB9_NOT1 = 2.7440
.param LRB1_NOT1 = 1.5503e-12
.param LRB2_NOT1 = 1.5081e-12
.param LRB3_NOT1 = 3.6223e-12
.param LRB4_NOT1 = 1.5503e-12
.param LRB5_NOT1 = 2.8924e-12
.param LRB6_NOT1 = 1.2792e-12
.param LRB7_NOT1 = 2.8086e-12
.param LRB8_NOT1 = 4.8448e-12
.param LRB9_NOT1 = 1.5503e-12
.param RD_NOT1 = 4
.param LRD_NOT1 = 2.0000e-12

B1_NOT1 1_NOT1 2_NOT1 jjmit_NOT1 area=B1_NOT1
B2_NOT1 4_NOT1 5_NOT1 jjmit_NOT1 area=B2_NOT1
B3_NOT1 7_NOT1 8_NOT1 jjmit_NOT1 area=B3_NOT1
B4_NOT1 13_NOT1 14_NOT1 jjmit_NOT1 area=B4_NOT1
B5_NOT1 17_NOT1 18_NOT1 jjmit_NOT1 area=B5_NOT1
B6_NOT1 10_NOT1 11_NOT1 jjmit_NOT1 area=B6_NOT1
B7_NOT1 20_NOT1 18_NOT1 jjmit_NOT1 area=B7_NOT1
B8_NOT1 18_NOT1 19_NOT1 jjmit_NOT1 area=B8_NOT1
B9_NOT1 21_NOT1 22_NOT1 jjmit_NOT1 area=B9_NOT1

IB1_NOT1 0 3_NOT1 pwl(0 0 5p IB1_NOT1)
IB2_NOT1 0 6_NOT1 pwl(0 0 5p IB2_NOT1)
IB3_NOT1 0 9_NOT1 pwl(0 0 5p IB3_NOT1)
IB4_NOT1 0 15_NOT1 pwl(0 0 5p IB4_NOT1)
IB5_NOT1 0 23_NOT1 pwl(0 0 5p IB5_NOT1)

LB1_NOT1 3_NOT1 1_NOT1 LB1_NOT1
LB2_NOT1 6_NOT1 4_NOT1 LB2_NOT1
LB3_NOT1 8_NOT1 9_NOT1 LB3_NOT1
LB4_NOT1 13_NOT1 15_NOT1 LB4_NOT1
LB5_NOT1 21_NOT1 23_NOT1 LB5_NOT1

L1_NOT1 a_NOT1 1_NOT1 2.062E-12
L2_NOT1 1_NOT1 4_NOT1 1.889E-12
L3_NOT1 4_NOT1 7_NOT1 2.72E-12
L4_NOT1 clk_NOT1 13_NOT1 2.057E-12
L5_NOT1 13_NOT1 16_NOT1 1.029E-12
L6_NOT1 16_NOT1 17_NOT1 1.241E-12
L7_NOT1 16_NOT1 12_NOT1 1.973E-12
L8_NOT1 10_NOT1 12_NOT1 1.003E-12
L9_NOT1 10_NOT1 8_NOT1 7.524E-12
L10_NOT1 8_NOT1 20_NOT1 1.234E-12
L11_NOT1 18_NOT1 21_NOT1 2.607E-12
L12_NOT1 21_NOT1 q_NOT1 2.062E-12

LP1_NOT1 2_NOT1 0 5.271E-13
LP2_NOT1 5_NOT1 0 5.237E-13
LP4_NOT1 14_NOT1 0 4.759E-13
LP6_NOT1 11_NOT1 0 5.021E-13
LP8_NOT1 19_NOT1 0 6.33E-13
LP9_NOT1 22_NOT1 0 4.749E-13

RB1_NOT1 1_NOT1 101_NOT1 RB1_NOT1
LRB1_NOT1 101_NOT1 0 LRB1_NOT1
RB2_NOT1 4_NOT1 104_NOT1 RB2_NOT1
LRB2_NOT1 104_NOT1 5_NOT1 LRB2_NOT1
RB3_NOT1 7_NOT1 107_NOT1 RB3_NOT1
LRB3_NOT1 107_NOT1 8_NOT1 LRB3_NOT1
RB4_NOT1 13_NOT1 113_NOT1 RB4_NOT1
LRB4_NOT1 113_NOT1 0 LRB4_NOT1
RB5_NOT1 17_NOT1 117_NOT1 RB5_NOT1
LRB5_NOT1 117_NOT1 18_NOT1 LRB5_NOT1
RB6_NOT1 10_NOT1 110_NOT1 RB6_NOT1
LRB6_NOT1 110_NOT1 0 LRB6_NOT1
RB7_NOT1 20_NOT1 120_NOT1 RB7_NOT1
LRB7_NOT1 120_NOT1 18_NOT1 LRB7_NOT1
RB8_NOT1 18_NOT1 118_NOT1 RB8_NOT1
LRB8_NOT1 118_NOT1 0 LRB8_NOT1
RB9_NOT1 21_NOT1 121_NOT1 RB9_NOT1
LRB9_NOT1 121_NOT1 0 LRB9_NOT1
LRD_NOT1 12_NOT1 112_NOT1 LRD_NOT1
RD_NOT1 112_NOT1 0 RD_NOT1
* .ends



*JTLNOT
LC_JTLNOT_1 CLKnn a_JTLNOT 0
LC_JTLNOT_2 CLK1nn q_JTLNOT 0

.model jjmit_JTLNOT jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLNOT = 2.0678e-15
.param B0_JTLNOT = 1
.param Ic0_JTLNOT = 1.0000e-04
.param IcRs_JTLNOT = 6.8599e-04
.param B0Rs_JTLNOT = 6.8599
.param Rsheet_JTLNOT = 2
.param Lsheet_JTLNOT = 1.1300e-12
.param LP_JTLNOT = 2.0000e-13
.param IC_JTLNOT = 2.5000
.param Lptl_JTLNOT = 2.0000e-12
.param LB_JTLNOT = 2.0000e-12
.param BiasCoef_JTLNOT = 0.7000
.param B1_JTLNOT = 2.5000
.param B2_JTLNOT = 2.5000
.param IB1_JTLNOT = 3.5000e-04
.param LB1_JTLNOT = 2.0000e-12
.param L1_JTLNOT = 2.0678e-12
.param L2_JTLNOT = 2.0678e-12
.param L3_JTLNOT = 2.0678e-12
.param L4_JTLNOT = 2.0678e-12
.param RB1_JTLNOT = 2.7440
.param RB2_JTLNOT = 2.7440
.param LRB1_JTLNOT = 1.7503e-12
.param LRB2_JTLNOT = 1.7503e-12
.param LP1_JTLNOT = 2.0000e-13
.param LP2_JTLNOT = 2.0000e-13

B1_JTLNOT 1_JTLNOT 2_JTLNOT jjmit_JTLNOT area=B1_JTLNOT
B2_JTLNOT 6_JTLNOT 7_JTLNOT jjmit_JTLNOT area=B2_JTLNOT
IB1_JTLNOT 0 5_JTLNOT pwl(0 0 5p IB1_JTLNOT)
L1_JTLNOT a_JTLNOT 1_JTLNOT 2.082E-12
L2_JTLNOT 1_JTLNOT 4_JTLNOT 2.06E-12
L3_JTLNOT 4_JTLNOT 6_JTLNOT 2.067E-12
L4_JTLNOT 6_JTLNOT q_JTLNOT 2.075E-12
LP1_JTLNOT 2_JTLNOT 0 4.998E-13
LP2_JTLNOT 7_JTLNOT 0 5.011E-13
LB1_JTLNOT 5_JTLNOT 4_JTLNOT LB1_JTLNOT
RB1_JTLNOT 1_JTLNOT 3_JTLNOT RB1_JTLNOT
RB2_JTLNOT 6_JTLNOT 8_JTLNOT RB2_JTLNOT
LRB1_JTLNOT 3_JTLNOT 0 LRB1_JTLNOT
LRB2_JTLNOT 8_JTLNOT 0 LRB2_JTLNOT
* .ends





.ends





