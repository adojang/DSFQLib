* A Generic Testbench for simulating Logic Gates
* Copyright (c) 2022-2024 Adriaan van Wijk, Stellenbosch University
*


.tran 0.25p 75p 0 0.025p

.param cval = 2.07m
.param ccval = 600u
.param Ic2 = 100u
.param Ic1 = 1.4 * Ic2
.param Ibx = 0.7 * Ic2

VsrcA B 0 pwl(0 0 30p 0 31p cval 32p 0 300p 0 301p cval 302p 0)

.model J2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=Ic2)

.model J1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=Ic1)

Ib 0 2 pwl(0 0 5p Ibx)


B2 1 2 J2
R2 1 22 2
L22 22 2 0.8p

B1 1 0 J1
R1 1 11 2
L11 11 0 0.8p

L1 A 1 2p
L2 2 B 2p

Rs A 0 2

.print p(1) p(2) p(B1) p(B2)


.end



* 2ps * 0.5 * 145
5ps * 0.5 * 164





*josim -o ./test.csv ./test.cir -V 1
*josim-plot.py ./test.csv -t stacked
