

.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_SFQDC_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include AW_mitll_DSFQ_OR.cir

.tran 0.025p 300p 0
.param cval= 600u
I_A0 0 xa pwl(0 0 100p 0 103p cval 105p 0 200p 0 203p cval 205p 0 300p 0 303p 0 305p 0) 
I_B0 0 xb pwl(0 0 105p 0 108p 0 110p 0 205p 0 208p cval 210p 0 315p 0 318p 0 320p 0)


XDCSFQA LSmitll_DCSFQ xa xa1 
XDCSFQB LSmitll_DCSFQ xb xb1
XDCSFQC LSmitll_DCSFQ xc xc1 
XDCSFQD LSmitll_DCSFQ xd xd1


XJTLA LSMITLL_JTL xa1 A
XJTLB LSMITLL_JTL xb1 B

XJTLC LSMITLL_JTL xc1 C
XJTLD LSMITLL_JTL xd1 D

* INSERT CELL HERE
XDUT DSFQ_OR A B q
* XDUT1 DSFQ_OR C D q

XLOAD LSMITLL_JTL q qq

Rsink qq 0 2
 .print i(L1.xdut) p(L2.XDUT) p(4.xdut) p(10.xdut) p(B6.xdut)  p(30.xdut) p(qq)
*  .print p(A) p(B) p(C) p(D) p(Q0) p(Q1) p(Q)
* .print p(q)

*110ps
*116.025ps
*Avg about 3ps
.end