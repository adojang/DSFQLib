.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_SFQDC_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include AW_mitll_DSFQ_OR.cir

.tran 0.015p 600p 0
.param cval= 600u
I_A0 0 xa pwl(0 0 100p 0 103p cval 105p 0 200p 0 203p cval 205p 0 300p 0 303p cval 305p 0 400p 0 403p cval 405p 0 500p 0 503p cval 505p 0) 
I_B0 0 xb pwl(0 0 110p 0 113p cval 115p 0 204p 0 207p 0 209p 0 306p 0 309p 0 311p 0 408p 0 411p 0 413p 0 510p 0 513p cval 515p 0)

XDCSFQA LSmitll_DCSFQ xa xa1 
XDCSFQB LSmitll_DCSFQ xb xb1

XJTLA LSMITLL_JTL xa1 A
XJTLB LSMITLL_JTL xb1 B

XDUT DSFQ_OR A B q

XLOAD LSMITLL_JTL q qq
Rsink qq 0 2

.print p(A) p(B) p(Q)
.end