* DSFQ Self clocked Multiplexor
* Author: Adriaan van Wijk
* Version: 1.0
* Last modification date: 21 June 2022
* Last modification by: Adriaan van Wijk
* This testbench uses cells from LS's library of RSFQ cells. This was the version that was tested for layout.

.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include cells\LSmitll_SPLIT_v2p1_optimized.cir
.include cells\LSmitll_NOT_v2p1_optimized.cir
.include AW_mitll_DSFQ_AND.cir
.include AW_mitll_DSFQ_OR.cir
.include AW_mitll_DSFQ_NOT.cir


.include newXOR.cir

.param cval=600u

I_a0 0 I_a0 pwl(0 0 100p 0 103p cval 105p 0        19p 0 110p 0 113p 0     300p 0 303p 0 305p 0     400p 0 403p 0 405p 0)
I_b0 0 I_b0 pwl(0 0 100p 0 103p 0 105p 0           140p 0 143p 0 145p 0       155p 0 158p cval 160p 0     300p 0 303p 0 305p 0        400p 0 403p 0 405p 0)
I_s0 0 I_s0 pwl(0 0 100p 0 103p cval 105p 0        110p 0 113p 0 115p 0        300p 0 303p 0 305p 0     400p 0 403p 0 405p 0)
I_m0 0 I_m0 pwl(0 0 100p 0 103p 0 105p 0        120p 0 123p cval 125p 0        300p 0 303p 0 305p 0     400p 0 403p 0 405p 0)

* A     0 0 1 1
* B     0 1 0 1
* AND1  0 0 0 1
* AND2  0 1 1 0
* Q     0 1 1 0

XSPLITtest LSmitll_SPLIT   S0      S1     S2

Xsrc_m0 LSmitll_DCSFQ i_m0 src_m0
*Feedback into SPLIT CELL
Xload_m0 LSMITLL_JTL src_m0 S2


RS1 S1 0 2

.tran 0.25p 300p 0 0.01p

Xsrc_a0 LSmitll_DCSFQ i_a0 src_a0
Xsrc_b0 LSmitll_DCSFQ i_b0 src_b0
Xsrc_s0 LSmitll_DCSFQ i_s0 src_s0

Xload_a0 LSMITLL_JTL src_a0 A0
Xload_b0 LSMITLL_JTL src_b0 B0
Xload_s0 LSMITLL_JTL src_s0 S0


XXOR DSFQ_XOR A0 B0 QQ

XLOAD LSMITLL_JTL QQ Qload
R_out Qload 0 2
XLOADS LSMITLL_JTL S0 Sout
R_REF Sout 0 2

* .print p(A0) p(B0) p(A11.xxor) p(B11.xxor) p(AND1.xxor) p(AND2.xxor) p(QQ) p(Sout)
* .print p(B4.XXOR) p(A4.XXOR) p(OR1.XXOR) p(OR2.XXOR) p(OR3.XXOR) p(B0) p(QQ) p(Sout)

.print p(S0) p(S1) p(S2)
 .print  p(A3.XXOR) p(src_b0) p(B0) p(B3.XXOR) p(AND1.XXOR) p(AND2.XXOR) p(B4.XXOR)



.end