.title KiCad schematic
LRB3 Net-_LRB3-Pad1_ Net-_B1-Pad1_ Inductor
RB4 Net-_B1-Pad1_ Net-_LRB4-Pad1_ Resistor
B6 Net-_B6-Pad1_ Net-_B2-Pad1_ jjmit
LRB4 Net-_LRB4-Pad1_ GND Inductor
RB5 Net-_B3-Pad2_ Net-_LRB5-Pad1_ Resistor
L3 Net-_B3-Pad2_ Net-_B8-Pad2_ Inductor
LRB5 Net-_LRB5-Pad1_ Net-_B2-Pad1_ Inductor
RB3 Net-_B3-Pad2_ Net-_LRB3-Pad1_ Resistor
I1 GND Net-_B3-Pad2_ pwl(0 0 100u)
RB6 Net-_B2-Pad1_ Net-_LRB6-Pad1_ Resistor
LP2 Net-_B6-Pad1_ GND Inductor
LRB6 Net-_LRB6-Pad1_ GND Inductor
B5 Net-_B2-Pad1_ Net-_B3-Pad2_ jjmit
RB9 Net-_B9-Pad2_ Net-_LRB9-Pad1_ Resistor
B9 Net-_B9-Pad1_ Net-_B9-Pad2_ jjmit
L4 Net-_B8-Pad2_ Net-_B7-Pad2_ Inductor
LRB7 Net-_LRB7-Pad1_ GND Inductor
LP3 Net-_B7-Pad1_ GND Inductor
LRB8 Net-_LRB8-Pad1_ Net-_B8-Pad1_ Inductor
RB8 Net-_B8-Pad2_ Net-_LRB8-Pad1_ Resistor
B8 Net-_B8-Pad1_ Net-_B8-Pad2_ jjmit
L5 Net-_B8-Pad1_ GND Inductor
L6 Net-_B8-Pad2_ Q Inductor
LP4 Net-_B9-Pad1_ GND Inductor
LRB9 Net-_LRB9-Pad1_ GND Inductor
R1 Net-_B7-Pad2_ Net-_B9-Pad2_ Resistor
B7 Net-_B7-Pad1_ Net-_B7-Pad2_ jjmit
RB7 Net-_B7-Pad2_ Net-_LRB7-Pad1_ Resistor
LP1 Net-_B4-Pad1_ GND Inductor
B4 Net-_B4-Pad1_ Net-_B1-Pad1_ jjmit
B1 Net-_B1-Pad1_ Net-_B1-Pad2_ jjmit
RB1 Net-_B1-Pad2_ Net-_LRB1-Pad1_ Resistor
LRB1 Net-_LRB1-Pad1_ Net-_B1-Pad1_ Inductor
RB2 Net-_B2-Pad2_ Net-_LRB2-Pad1_ Resistor
B2 Net-_B2-Pad1_ Net-_B2-Pad2_ jjmit
LRB2 Net-_LRB2-Pad1_ Net-_B2-Pad1_ Inductor
L1 A Net-_B1-Pad2_ Inductor
L2 B Net-_B2-Pad2_ Inductor
B3 Net-_B1-Pad1_ Net-_B3-Pad2_ jjmit
.end
