* Author: Adriaan van Wijk
* Version: 1.2
* Last modification date: 28 March 2022
* Last modification by: Adriaan van Wijk
* Based on the design by Rylov [2019]

* Copyright (c) 2022 Adriaan van Wijk, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Adriaan van Wijk, 21786275@sun.ac.za

*$Ports    A B q
.subckt DSFQ_AND A B q

.param Ibias=70u
.param main=0.84
.param secondary=0.60
.param third=1.68

.param L1=8p
.param L2=8p
.param Lout=2p

* The throughput for this logic cell is approximately 5ps with zero skew applied.
* The skew tolerance can be adjusted using the following formula:
* RHold = a * (16.666 * t_hold)^b
* Where a = 3.572e-10
* and   b = -1.023

.param RHold = 3.597
.param RS = RHold
.param RD = RHold

*The precalculated values for the parasitic inductances and resistances
.param RBA=11.4332
.param LBA=6.4597p
.param RBB=8.1666
.param LBB=4.6141p
.param RBC=4.0833
.param LBC=2.3071p

L1 A 1 L1
L2 B 4 L2

RD1 1 2 RD
RD2 4 5 RD
BD1 2 C jjmit area=secondary
RDp1 2 14 RBA
Ld1 14 C LBA

BD2 5 C jjmit area=secondary
RDp2 5 15 RBA
Ld2 15 C LBA
RS1 1 C RS
RS2 4 C RS

B1 1 C jjmit area=main
Rb1 1 10 RBB
Lb1 10 C LBB

B2 4 C jjmit area=main
Rb2 4 11 RBB
Lb2 11 C LBB

B3 C 0 jjmit area=third
Rb3 C 13 RBC
Lb3 13 0 LBC

Ibias 0 C dc Ibias
Lout q C Lout
.ends