.title KiCad schematic
I1 GND Net-_B1-Pad1_ pwl(0 0 100u)
B4 Net-_B2-Pad1_ Net-_B1-Pad1_ jjmit
LRB4 Net-_LRB4-Pad1_ Net-_B2-Pad1_ Inductor
RB4 Net-_B1-Pad1_ Net-_LRB4-Pad1_ Resistor
LRB3 Net-_LRB3-Pad1_ Net-_B1-Pad1_ Inductor
RB3 Net-_B3-Pad2_ Net-_LRB3-Pad1_ Resistor
B3 Net-_B1-Pad1_ Net-_B3-Pad2_ jjmit
L3 Net-_B1-Pad1_ Out Inductor
B5 Net-_B5-Pad1_ Net-_B1-Pad1_ jjmit
RB5 Net-_B1-Pad1_ Net-_LRB5-Pad1_ Resistor
LRB5 Net-_LRB5-Pad1_ GND Inductor
LP1 Net-_B5-Pad1_ GND Inductor
L2 B Net-_B2-Pad2_ Inductor
L1 A Net-_B1-Pad2_ Inductor
R1 Net-_B3-Pad2_ Net-_B1-Pad2_ Resistor
RB1 Net-_B1-Pad2_ Net-_LRB1-Pad1_ Resistor
LRB1 Net-_LRB1-Pad1_ Net-_B1-Pad1_ Inductor
R4 Net-_B2-Pad2_ Net-_B2-Pad1_ Resistor
B2 Net-_B2-Pad1_ Net-_B2-Pad2_ jjmit
R3 Net-_B1-Pad2_ Net-_B1-Pad1_ Resistor
B1 Net-_B1-Pad1_ Net-_B1-Pad2_ jjmit
RB2 Net-_B2-Pad2_ Net-_LRB2-Pad1_ Resistor
R2 Net-_B1-Pad1_ Net-_B2-Pad2_ Resistor
LRB2 Net-_LRB2-Pad1_ Net-_B2-Pad1_ Inductor
.end
