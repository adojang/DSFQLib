.title KiCad schematic
L7 /13 /16 Inductor
L6 /12 /13 Inductor
B7 /8 /12 jjmit
LP3 /8 GND Inductor
B9 /15 /17 jjmit
LP5 /15 GND Inductor
I2 GND /4 pwl(0 0 5p REF)
B6 /12 /4 jjmit
LP4 /14 GND Inductor
B8 /14 /13 jjmit
I3 GND /16 pwl(0 0 5p REF)
L8 /16 /17 Inductor
L9 /17 Q Inductor
L4 /10 /11 Inductor
L5 A /44 Inductor
B2 /6 /5 jjmit
LP1 /6 GND Inductor
L3 /9 /10 Inductor
I1 GND /9 pwl(0 0 5p REF)
B4 /12 /11 jjmit
B5 /4 /44 jjmit
L2 /5 /9 Inductor
LP2 /7 GND Inductor
B3 /7 /10 jjmit
B1 /5 /55 jjmit
L1 CLK /55 Inductor
.end
