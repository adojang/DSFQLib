.subckt SHUNT a b q
.param l1       =                3.09037291e-12
.param l3       =                2.03058886e-12
.param r1       =                7.04349127e-01
.param r3       =                1.34323634e+00
.param i1    =                40u

.param l2       =         l1
.param r2       =         r1
.param r4       =         r3

*Static Parameters
.param b1       =         5.16417451e-01
.param b2       =         b1
.param b3       =         3.3e-01
.param b4       =         b3
.param b5       =         1.05188201e+00

.param rb1      =         12.92859137e+00
.param rb2      =         12.92013085e+00
.param rb3      =         19.98871344e+00
.param rb4      =         19.98963516e+00
.param rb5      =         6.566007373e+00

.param lrb1     =         3.94321337e-13
.param lrb2     =         5.33421859e-13
.param lrb3     =         1.39314087e-12
.param lrb4     =         1.41001012e-12
.param lrb5     =         1.19776828e-12
.param lp1      =         8.25215763e-13

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
* Annotated .cir file from KiCad
b1   	30   	10   	 jjmit area=b1
b2   	30   	20   	 jjmit area=b2
b3   	30   	12   	 jjmit area=b3
b4   	30   	22   	 jjmit area=b4
b5   	31   	30   	 jjmit area=b5
i1   	0   	30   	pwl(0   	0   	5p   	i1)
l1   	a   	10   	 l1
l2   	b   	20   	 l2
l3   	30   	q   	 l3
lp1   	31   	0   	 lp1
lrb1   	11   	30   	 lrb1
lrb2   	21   	30   	 lrb2
lrb3   	net-_lrb3-pad1_   	30   	 lrb3
lrb4   	net-_lrb4-pad1_   	30   	 lrb4
lrb5   	32   	0   	 lrb5
r1   	10   	30   	 r1
r2   	20   	30   	 r2
r3   	12   	10   	 r3
r4   	22   	20   	 r4
rb1   	10   	11   	 rb1
rb2   	20   	21   	 rb2
rb3   	12   	net-_lrb3-pad1_   	 rb3
rb4   	22   	net-_lrb4-pad1_   	 rb4
rb5   	30   	32   	 rb5
.ends