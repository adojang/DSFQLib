
.subckt DSFQ_XOR A0 B0 QQ
*OPTIMIZED TESTBENCH 2.71 Margin on B9_NOT_NOT.



* XXOR DSFQ_XOR A0 B0 QQ
LXOR1 A0 A 0
LXOR2 B0 B 0
LXOR3 QQ Q 0


*THIS SUBCIRCUIT WAS FLATTENED. THE AND GATE HAS A SLIGHTLY SMALLER OUTPUT INDUCTANCE THAN IS TYPICAL, WHICH MAY CHANGE THE NORMAL MARGINS.


* .SUBCKT DSFQ_XOR A B Q

* XSPLITA LSMITLL_SPLITO A A1 A2
* XSPLITB LSMITLL_SPLITO B B1 B2

* XJTL1 LSMITLL_JTLI A1 A11
* XJTL2 LSMITLL_JTLI B1 B11
* XJTL3 LSMITLL_JTLI OR1 OR2
* XJTL4 LSMITLL_JTLI OR2 OR3

* XNAND1  DSFQ_ANDO    A1     B1   AND1
* XNAND2  DSFQ_NOTO    AND1   A11   B11   AND2
* XOR     DSFQ_ORI     A1     B2   OR1
* XAND    DSFQ_ANDO    AND2   OR3  Q

*LIBRARIES SO THE CIRCUIT CAN RUN BY ITSELF WITHOUT REQUIRING THE USER TO ADD THEM.
*LIBRARIES INCLUDED: DSFQ_AND DSFQ_OR LSMITLL_JTL, LSMITLL_SPLIT, LSMITLL_NOT DSFQ_NOT, 


*****JTL CELLS ***********************************************
*JTLA1
LC_JTLA1_1 A1 A_JTLA1 0
LC_JTLA1_2 A11 Q_JTLA1 0

.MODEL JJMIT_JTLA1 JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.PARAM PHI0_JTLA1 = 2.0678E-15
.PARAM B0_JTLA1 = 1
.PARAM IC0_JTLA1 = 1.0000E-04
.PARAM ICRS_JTLA1 = 6.8599E-04
.PARAM B0RS_JTLA1 = 6.8599
.PARAM RSHEET_JTLA1 = 2
.PARAM LSHEET_JTLA1 = 1.1300E-12
.PARAM LP_JTLA1 = 2.0000E-13
.PARAM IC_JTLA1 = 2.5000
.PARAM LPTL_JTLA1 = 2.0000E-12
.PARAM LB_JTLA1 = 2.0000E-12
.PARAM BIASCOEF_JTLA1 = 0.7000
.PARAM B1_JTLA1=2.516413e+00
.PARAM B2_JTLA1 = 2.5000
.PARAM IB1_JTLA1 = 3.5000E-04
.PARAM LB1_JTLA1 = 2.0000E-12
.PARAM L1_JTLA1 = 2.0678E-12
.PARAM L2_JTLA1 = 2.0678E-12
.PARAM L3_JTLA1 = 2.0678E-12
.PARAM L4_JTLA1 = 2.0678E-12
.PARAM RB1_JTLA1 = 2.7440
.PARAM RB2_JTLA1 = 2.7440
.PARAM LRB1_JTLA1 = 1.7503E-12
.PARAM LRB2_JTLA1 = 1.7503E-12
.PARAM LP1_JTLA1 = 2.0000E-13
.PARAM LP2_JTLA1 = 2.0000E-13

B1_JTLA1 1_JTLA1 2_JTLA1 JJMIT_JTLA1 AREA=B1_JTLA1
B2_JTLA1 6_JTLA1 7_JTLA1 JJMIT_JTLA1 AREA=B2_JTLA1
IB1_JTLA1 0 5_JTLA1 PWL(0 0 5P IB1_JTLA1)
L1_JTLA1 A_JTLA1 1_JTLA1 2.082E-12
L2_JTLA1 1_JTLA1 4_JTLA1 2.06E-12
L3_JTLA1 4_JTLA1 6_JTLA1 2.067E-12
L4_JTLA1 6_JTLA1 Q_JTLA1 2.075E-12
LP1_JTLA1 2_JTLA1 0 4.998E-13
LP2_JTLA1 7_JTLA1 0 5.011E-13
LB1_JTLA1 5_JTLA1 4_JTLA1 LB1_JTLA1
RB1_JTLA1 1_JTLA1 3_JTLA1 RB1_JTLA1
RB2_JTLA1 6_JTLA1 8_JTLA1 RB2_JTLA1
LRB1_JTLA1 3_JTLA1 0 LRB1_JTLA1
LRB2_JTLA1 8_JTLA1 0 LRB2_JTLA1

*JTLA2
LC_JTLA2_1 B1 A_JTLA2 0
LC_JTLA2_2 B11 Q_JTLA2 0

.MODEL JJMIT_JTLA2 JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.PARAM PHI0_JTLA2 = 2.0678E-15
.PARAM B0_JTLA2 = 1
.PARAM IC0_JTLA2 = 1.0000E-04
.PARAM ICRS_JTLA2 = 6.8599E-04
.PARAM B0RS_JTLA2 = 6.8599
.PARAM RSHEET_JTLA2 = 2
.PARAM LSHEET_JTLA2 = 1.1300E-12
.PARAM LP_JTLA2 = 2.0000E-13
.PARAM IC_JTLA2 = 2.5000
.PARAM LPTL_JTLA2 = 2.0000E-12
.PARAM LB_JTLA2 = 2.0000E-12
.PARAM BIASCOEF_JTLA2 = 0.7000
.PARAM B1_JTLA2 = 2.5000
.PARAM B2_JTLA2 = 2.5000
.PARAM IB1_JTLA2 = 3.5000E-04
.PARAM LB1_JTLA2 = 2.0000E-12
.PARAM L1_JTLA2 = 2.0678E-12
.PARAM L2_JTLA2 = 2.0678E-12
.PARAM L3_JTLA2 = 2.0678E-12
.PARAM L4_JTLA2 = 2.0678E-12
.PARAM RB1_JTLA2 = 2.7440
.PARAM RB2_JTLA2 = 2.7440
.PARAM LRB1_JTLA2 = 1.7503E-12
.PARAM LRB2_JTLA2 = 1.7503E-12
.PARAM LP1_JTLA2 = 2.0000E-13
.PARAM LP2_JTLA2 = 2.0000E-13

B1_JTLA2 1_JTLA2 2_JTLA2 JJMIT_JTLA2 AREA=B1_JTLA2
B2_JTLA2 6_JTLA2 7_JTLA2 JJMIT_JTLA2 AREA=B2_JTLA2
IB1_JTLA2 0 5_JTLA2 PWL(0 0 5P IB1_JTLA2)
L1_JTLA2 A_JTLA2 1_JTLA2 2.082E-12
L2_JTLA2 1_JTLA2 4_JTLA2 2.06E-12
L3_JTLA2 4_JTLA2 6_JTLA2 2.067E-12
L4_JTLA2 6_JTLA2 Q_JTLA2 2.075E-12
LP1_JTLA2 2_JTLA2 0 4.998E-13
LP2_JTLA2 7_JTLA2 0 5.011E-13
LB1_JTLA2 5_JTLA2 4_JTLA2 LB1_JTLA2
RB1_JTLA2 1_JTLA2 3_JTLA2 RB1_JTLA2
RB2_JTLA2 6_JTLA2 8_JTLA2 RB2_JTLA2
LRB1_JTLA2 3_JTLA2 0 LRB1_JTLA2
LRB2_JTLA2 8_JTLA2 0 LRB2_JTLA2

*JTLA3
LC_JTLA3_1 OR1 A_JTLA3 0
LC_JTLA3_2 OR2 Q_JTLA3 0

.MODEL JJMIT_JTLA3 JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.PARAM PHI0_JTLA3 = 2.0678E-15
.PARAM B0_JTLA3 = 1
.PARAM IC0_JTLA3 = 1.0000E-04
.PARAM ICRS_JTLA3 = 6.8599E-04
.PARAM B0RS_JTLA3 = 6.8599
.PARAM RSHEET_JTLA3 = 2
.PARAM LSHEET_JTLA3 = 1.1300E-12
.PARAM LP_JTLA3 = 2.0000E-13
.PARAM IC_JTLA3 = 2.5000
.PARAM LPTL_JTLA3 = 2.0000E-12
.PARAM LB_JTLA3 = 2.0000E-12
.PARAM BIASCOEF_JTLA3 = 0.7000
.PARAM B1_JTLA3 = 2.5000
.PARAM B2_JTLA3 = 2.5000
.PARAM IB1_JTLA3 = 3.5000E-04
.PARAM LB1_JTLA3 = 2.0000E-12
.PARAM L1_JTLA3 = 2.0678E-12
.PARAM L2_JTLA3 = 2.0678E-12
.PARAM L3_JTLA3 = 2.0678E-12
.PARAM L4_JTLA3 = 2.0678E-12
.PARAM RB1_JTLA3 = 2.7440
.PARAM RB2_JTLA3 = 2.7440
.PARAM LRB1_JTLA3 = 1.7503E-12
.PARAM LRB2_JTLA3 = 1.7503E-12
.PARAM LP1_JTLA3 = 2.0000E-13
.PARAM LP2_JTLA3 = 2.0000E-13

B1_JTLA3 1_JTLA3 2_JTLA3 JJMIT_JTLA3 AREA=B1_JTLA3
B2_JTLA3 6_JTLA3 7_JTLA3 JJMIT_JTLA3 AREA=B2_JTLA3
IB1_JTLA3 0 5_JTLA3 PWL(0 0 5P IB1_JTLA3)
L1_JTLA3 A_JTLA3 1_JTLA3 2.082E-12
L2_JTLA3 1_JTLA3 4_JTLA3 2.06E-12
L3_JTLA3 4_JTLA3 6_JTLA3 2.067E-12
L4_JTLA3 6_JTLA3 Q_JTLA3 2.075E-12
LP1_JTLA3 2_JTLA3 0 4.998E-13
LP2_JTLA3 7_JTLA3 0 5.011E-13
LB1_JTLA3 5_JTLA3 4_JTLA3 LB1_JTLA3
RB1_JTLA3 1_JTLA3 3_JTLA3 RB1_JTLA3
RB2_JTLA3 6_JTLA3 8_JTLA3 RB2_JTLA3
LRB1_JTLA3 3_JTLA3 0 LRB1_JTLA3
LRB2_JTLA3 8_JTLA3 0 LRB2_JTLA3

*JTLA4
LC_JTLA4_1 OR2 A_JTLA4 0
LC_JTLA4_2 OR3 Q_JTLA4 0

.MODEL JJMIT_JTLA4 JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.PARAM PHI0_JTLA4 = 2.0678E-15
.PARAM B0_JTLA4 = 1
.PARAM IC0_JTLA4 = 1.0000E-04
.PARAM ICRS_JTLA4 = 6.8599E-04
.PARAM B0RS_JTLA4 = 6.8599
.PARAM RSHEET_JTLA4 = 2
.PARAM LSHEET_JTLA4 = 1.1300E-12
.PARAM LP_JTLA4 = 2.0000E-13
.PARAM IC_JTLA4 = 2.5000
.PARAM LPTL_JTLA4 = 2.0000E-12
.PARAM LB_JTLA4 = 2.0000E-12
.PARAM BIASCOEF_JTLA4 = 0.7000
.PARAM B1_JTLA4 = 2.5000
.PARAM B2_JTLA4 = 2.5000
.PARAM IB1_JTLA4 = 3.5000E-04
.PARAM LB1_JTLA4 = 2.0000E-12
.PARAM L1_JTLA4 = 2.0678E-12
.PARAM L2_JTLA4 = 2.0678E-12
.PARAM L3_JTLA4 = 2.0678E-12
.PARAM L4_JTLA4 = 2.0678E-12
.PARAM RB1_JTLA4 = 2.7440
.PARAM RB2_JTLA4 = 2.7440
.PARAM LRB1_JTLA4 = 1.7503E-12
.PARAM LRB2_JTLA4 = 1.7503E-12
.PARAM LP1_JTLA4 = 2.0000E-13
.PARAM LP2_JTLA4 = 2.0000E-13

B1_JTLA4 1_JTLA4 2_JTLA4 JJMIT_JTLA4 AREA=B1_JTLA4
B2_JTLA4 6_JTLA4 7_JTLA4 JJMIT_JTLA4 AREA=B2_JTLA4
IB1_JTLA4 0 5_JTLA4 PWL(0 0 5P IB1_JTLA4)
L1_JTLA4 A_JTLA4 1_JTLA4 2.082E-12
L2_JTLA4 1_JTLA4 4_JTLA4 2.06E-12
L3_JTLA4 4_JTLA4 6_JTLA4 2.067E-12
L4_JTLA4 6_JTLA4 Q_JTLA4 2.075E-12
LP1_JTLA4 2_JTLA4 0 4.998E-13
LP2_JTLA4 7_JTLA4 0 5.011E-13
LB1_JTLA4 5_JTLA4 4_JTLA4 LB1_JTLA4
RB1_JTLA4 1_JTLA4 3_JTLA4 RB1_JTLA4
RB2_JTLA4 6_JTLA4 8_JTLA4 RB2_JTLA4
LRB1_JTLA4 3_JTLA4 0 LRB1_JTLA4
LRB2_JTLA4 8_JTLA4 0 LRB2_JTLA4




*AND1

LC_AND1_1 A1 A_AND1 0
LC_AND1_2 B1 B_AND1 0
LC_AND1_3 AND1 Q_AND1 0

.PARAM B1_AND1 = 1.39878486E+00
.PARAM BD1_AND1 = 1.38855937E+00
.PARAM L1_AND1 = 1.64204687E-12
.PARAM RD1_AND1 = 6.00718616E-01
.PARAM I1_AND1 = 1.54457273E-05
.PARAM B3_AND1 = 1.51517089E+00
*THIS LINE WAS EDITED TO MAKE THE SIMULATION WORK
*THIS MIGHT CHANGE THE WHOLE MARGINS OF THE FILE. NEED TO CHECK IF AND IS STILL OKAY WITH THIS.
.PARAM L3_AND1 = 4.24567618E-13
.PARAM RH1_AND1 = 4.76237371E+00
.PARAM LDP1_AND1 = 1E-12
.PARAM B2_AND1 = B1_AND1
.PARAM BD2_AND1 = BD1_AND1
.PARAM L2_AND1 = L1_AND1
.PARAM LDP2_AND1 = LDP1_AND1
.PARAM RD2_AND1 = RD1_AND1
.PARAM LP1_AND1 = 0.2E-12
.PARAM LHP1_AND1 = 1E-12
.PARAM LHP2_AND1 = LHP1_AND1
.PARAM RH2_AND1 = RH1_AND1

.MODEL JJMIT_AND1 JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)

B1_AND1 30_AND1 10_AND1 JJMIT_AND1 AREA=B1_AND1
B2_AND1 30_AND1 20_AND1 JJMIT_AND1 AREA=B2_AND1
B3_AND1 31_AND1 30_AND1 JJMIT_AND1 AREA=B3_AND1
BD1_AND1 30_AND1 12_AND1 JJMIT_AND1 AREA=BD1_AND1
BD2_AND1 30_AND1 22_AND1 JJMIT_AND1 AREA=BD2_AND1
I1_AND1 0 30_AND1 PWL(0 0 5P I1_AND1)
L1_AND1 A_AND1 10_AND1 L1_AND1
L2_AND1 B_AND1 20_AND1 L2_AND1
L3_AND1 30_AND1 Q_AND1 L3_AND1
LDP1_AND1 11_AND1 12_AND1 LDP1_AND1
LDP2_AND1 21_AND1 22_AND1 LDP2_AND1
LHP1_AND1 13_AND1 30_AND1 LHP1_AND1
LHP2_AND1 23_AND1 30_AND1 LHP2_AND1
LP1_AND1 31_AND1 0 LP1_AND1
RD1_AND1 11_AND1 10_AND1 RD1_AND1
RD2_AND1 21_AND1 20_AND1 RD2_AND1
RH1_AND1 13_AND1 10_AND1 RH1_AND1
RH2_AND1 23_AND1 20_AND1 RH2_AND1


*AND2

LC_AND2_1 AND2 A_AND2 0
LC_AND2_2 OR3 B_AND2 0
LC_AND2_3 Q Q_AND2 0

.PARAM B1_AND2 = 1.39878486E+00
.PARAM BD1_AND2 = 1.38855937E+00
.PARAM L1_AND2 = 1.64204687E-12
.PARAM RD1_AND2 = 6.00718616E-01
.PARAM I1_AND2 = 1.54457273E-05
.PARAM B3_AND2=1.484143e+00
*THIS LINE WAS EDITED TO MAKE THE SIMULATION WORK
*THIS MIGHT CHANGE THE WHOLE MARGINS OF THE FILE. NEED TO CHECK IF AND IS STILL OKAY WITH THIS.
.PARAM L3_AND2 = 4.24567618E-13
.PARAM RH1_AND2 = 4.76237371E+00
.PARAM LDP1_AND2 = 1E-12
.PARAM B2_AND2 = B1_AND2
.PARAM BD2_AND2 = BD1_AND2
.PARAM L2_AND2 = L1_AND2
.PARAM LDP2_AND2 = LDP1_AND2
.PARAM RD2_AND2 = RD1_AND2
.PARAM LP1_AND2 = 0.2E-12
.PARAM LHP1_AND2 = 1E-12
.PARAM LHP2_AND2 = LHP1_AND2
.PARAM RH2_AND2 = RH1_AND2

.MODEL JJMIT_AND2 JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)

B1_AND2 30_AND2 10_AND2 JJMIT_AND2 AREA=B1_AND2
B2_AND2 30_AND2 20_AND2 JJMIT_AND2 AREA=B2_AND2
B3_AND2 31_AND2 30_AND2 JJMIT_AND2 AREA=B3_AND2
BD1_AND2 30_AND2 12_AND2 JJMIT_AND2 AREA=BD1_AND2
BD2_AND2 30_AND2 22_AND2 JJMIT_AND2 AREA=BD2_AND2
I1_AND2 0 30_AND2 PWL(0 0 5P I1_AND2)
L1_AND2 A_AND2 10_AND2 L1_AND2
L2_AND2 B_AND2 20_AND2 L2_AND2
L3_AND2 30_AND2 Q_AND2 L3_AND2
LDP1_AND2 11_AND2 12_AND2 LDP1_AND2
LDP2_AND2 21_AND2 22_AND2 LDP2_AND2
LHP1_AND2 13_AND2 30_AND2 LHP1_AND2
LHP2_AND2 23_AND2 30_AND2 LHP2_AND2
LP1_AND2 31_AND2 0 LP1_AND2
RD1_AND2 11_AND2 10_AND2 RD1_AND2
RD2_AND2 21_AND2 20_AND2 RD2_AND2
RH1_AND2 13_AND2 10_AND2 RH1_AND2
RH2_AND2 23_AND2 20_AND2 RH2_AND2




* XOR     DSFQ_ORI     A1     B2   OR1

LC_OR1_1 A1 A_OR1 0
LC_OR1_2 B2 B_OR1 0
LC_OR1_3 OR1 Q_OR1 0

* .SUBCKT DSFQ_OR1 A_OR1 B_OR1 Q_OR1
.MODEL JJMIT_OR1 JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
*CONFLUENCE BUFFER A
.PARAM L1_OR1 = 2E-12
.PARAM B1_OR1 = 1.37211310E+00
.PARAM B3_OR1 = 2.77209629E+00
.PARAM B4_OR1 = 3.78734058E-01

* AND GATE LOOP
.PARAM L4_OR1 = 1.22182342E-12
.PARAM B7_OR1 = 1.19265113E+00
.PARAM B9_OR1 = 5.40924075E-01
.PARAM L7_OR1 = 1.62539785E-13
.PARAM R1_OR1 = 1.09745275E+01
.PARAM R2_OR1 = 5.58089917E-01
.PARAM L5_OR1 = 5.61756493E-13

* OUTPUT STAGE
.PARAM B8_OR1 = 7.09413113E-01
.PARAM I1_OR1 = 3.23631555E-04
.PARAM L3_OR1 = 2E-12
.PARAM L6_OR1 = 3.06315548E-12

*CONFLUENCE BUFFER B
.PARAM L2_OR1 = L1_OR1
.PARAM B2_OR1 = B1_OR1
.PARAM B5_OR1 = B3_OR1
.PARAM B6_OR1 = B4_OR1

*PARASITICS
.PARAM LP1_OR1 = 0.2E-12
.PARAM LP2_OR1 = 0.2E-12
.PARAM LP3_OR1 = 0.2E-12
.PARAM LP4_OR1 = 0.2E-12

* BACK ANNOTATED .CIR FILE FROM KICAD
B1_OR1 3_OR1 1_OR1 JJMIT_OR1 AREA=B1_OR1
B2_OR1 4_OR1 2_OR1 JJMIT_OR1 AREA=B2_OR1
B3_OR1 3_OR1 10_OR1 JJMIT_OR1 AREA=B3_OR1
B4_OR1 5_OR1 3_OR1 JJMIT_OR1 AREA=B4_OR1
B5_OR1 4_OR1 10_OR1 JJMIT_OR1 AREA=B5_OR1
B6_OR1 6_OR1 4_OR1 JJMIT_OR1 AREA=B6_OR1
B7_OR1 24_OR1 20_OR1 JJMIT_OR1 AREA=B7_OR1
B8_OR1 30_OR1 31_OR1 JJMIT_OR1 AREA=B8_OR1
B9_OR1 24_OR1 23_OR1 JJMIT_OR1 AREA=B9_OR1
I1_OR1 0 10_OR1 PWL(0 0 5P I1_OR1)
L1_OR1 A_OR1 1_OR1 L1_OR1
L2_OR1 B_OR1 2_OR1 L2_OR1
L3_OR1 10_OR1 30_OR1 L3_OR1
L4_OR1 30_OR1 20_OR1 L4_OR1
L5_OR1 21_OR1 24_OR1 L5_OR1
L6_OR1 30_OR1 Q_OR1 L6_OR1
L7_OR1 22_OR1 23_OR1 L7_OR1
LP1_OR1 5_OR1 0 LP1_OR1
LP2_OR1 6_OR1 0 LP2_OR1
LP3_OR1 24_OR1 0 LP3_OR1
LP4_OR1 31_OR1 0 LP4_OR1
R1_OR1 21_OR1 20_OR1 R1_OR1
R2_OR1 22_OR1 20_OR1 R2_OR1




* XNAND2  DSFQ_NOTO    AND1   A11   B11   AND2

LC_NOT_1 ANNN AND1 0
LC_NOT_2 BNNN A11 0
LC_NOT_3 CNNN B11 0
LC_NOT_4 QNNN AND2 0

*************** NEW NOT GATE
* .SUBCKT DSFQ_NOTO A B C Q
* .MODEL JJMIT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
*A IS INVERTING INPUT.
*B AND C ARE INPUTS FOR THE OR GATE.
*Q IS OUTPUT.

* XDSFQ_OR DSFQ_ORI B C CLKD
* XJTLCLK LSMITLL_JTLI CLKD CLK
* XNOTLS LSMITLL_NOTI A CLK Q

*NNOT

LC_NOT_NOT_1 ANNN A_NOT_NOT 0
LC_NOT_NOT_2 CLK CLK_NOT_NOT 0
LC_NOT_NOT_3 QNNN Q_NOT_NOT 0
* .SUBCKT LSMITLL_NOTI_NOT_NOT A_NOT_NOT CLK_NOT_NOT Q_NOT_NOT
.MODEL JJMIT_NOT_NOT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.PARAM PHI0_NOT_NOT = 2.0678E-15
.PARAM B0_NOT_NOT = 1
.PARAM IC0_NOT_NOT = 1.0000E-04
.PARAM ICRS_NOT_NOT = 6.8599E-04
.PARAM B0RS_NOT_NOT = 6.8599
.PARAM RSHEET_NOT_NOT = 2
.PARAM LSHEET_NOT_NOT = 1.1300E-12
.PARAM LP_NOT_NOT = 2.0000E-13
.PARAM IC_NOT_NOT = 2.5000
.PARAM LB_NOT_NOT = 2.0000E-12
.PARAM BIASCOEF_NOT_NOT = 0.7000
.PARAM B1_NOT_NOT = 2.5000
.PARAM B2_NOT_NOT = 2.5700
.PARAM B3_NOT_NOT = 1.0700
.PARAM B4_NOT_NOT = 2.5000
.PARAM B5_NOT_NOT=1.160533e+00
.PARAM B6_NOT_NOT = 3.0300
.PARAM B7_NOT_NOT = 1.3800
.PARAM B8_NOT_NOT=8.437228e-01
.PARAM B9_NOT_NOT=2.667062e+00
.PARAM IB1_NOT_NOT = 1.7500E-04
.PARAM IB2_NOT_NOT = 8.7000E-05
.PARAM IB3_NOT_NOT=2.509517e-04
.PARAM IB4_NOT_NOT = 1.7500E-04
.PARAM IB5_NOT_NOT = 1.7500E-04
.PARAM LB1_NOT_NOT = 2.0000E-12
.PARAM LB2_NOT_NOT = 2.0000E-12
.PARAM LB3_NOT_NOT = 2.0000E-12
.PARAM LB4_NOT_NOT = 2.0000E-12
.PARAM LB5_NOT_NOT = 2.0000E-12
.PARAM RB1_NOT_NOT = 2.7440
.PARAM RB2_NOT_NOT = 2.6692
.PARAM RB3_NOT_NOT = 6.4111
.PARAM RB4_NOT_NOT = 2.7440
.PARAM RB5_NOT_NOT = 5.1193
.PARAM RB6_NOT_NOT = 2.2640
.PARAM RB7_NOT_NOT = 4.9709
.PARAM RB8_NOT_NOT = 8.5749
.PARAM RB9_NOT_NOT = 2.7440
.PARAM LRB1_NOT_NOT = 1.5503E-12
.PARAM LRB2_NOT_NOT = 1.5081E-12
.PARAM LRB3_NOT_NOT = 3.6223E-12
.PARAM LRB4_NOT_NOT = 1.5503E-12
.PARAM LRB5_NOT_NOT = 2.8924E-12
.PARAM LRB6_NOT_NOT = 1.2792E-12
.PARAM LRB7_NOT_NOT = 2.8086E-12
.PARAM LRB8_NOT_NOT = 4.8448E-12
.PARAM LRB9_NOT_NOT = 1.5503E-12
.PARAM RD_NOT_NOT = 4
.PARAM LRD_NOT_NOT = 2.0000E-12

B1_NOT_NOT 1_NOT_NOT 2_NOT_NOT JJMIT_NOT_NOT AREA=B1_NOT_NOT
B2_NOT_NOT 4_NOT_NOT 5_NOT_NOT JJMIT_NOT_NOT AREA=B2_NOT_NOT
B3_NOT_NOT 7_NOT_NOT 8_NOT_NOT JJMIT_NOT_NOT AREA=B3_NOT_NOT
B4_NOT_NOT 13_NOT_NOT 14_NOT_NOT JJMIT_NOT_NOT AREA=B4_NOT_NOT
B5_NOT_NOT 17_NOT_NOT 18_NOT_NOT JJMIT_NOT_NOT AREA=B5_NOT_NOT
B6_NOT_NOT 10_NOT_NOT 11_NOT_NOT JJMIT_NOT_NOT AREA=B6_NOT_NOT
B7_NOT_NOT 20_NOT_NOT 18_NOT_NOT JJMIT_NOT_NOT AREA=B7_NOT_NOT
B8_NOT_NOT 18_NOT_NOT 19_NOT_NOT JJMIT_NOT_NOT AREA=B8_NOT_NOT
B9_NOT_NOT 21_NOT_NOT 22_NOT_NOT JJMIT_NOT_NOT AREA=B9_NOT_NOT

IB1_NOT_NOT 0 3_NOT_NOT PWL(0 0 5P IB1_NOT_NOT)
IB2_NOT_NOT 0 6_NOT_NOT PWL(0 0 5P IB2_NOT_NOT)
IB3_NOT_NOT 0 9_NOT_NOT PWL(0 0 5P IB3_NOT_NOT)
IB4_NOT_NOT 0 15_NOT_NOT PWL(0 0 5P IB4_NOT_NOT)
IB5_NOT_NOT 0 23_NOT_NOT PWL(0 0 5P IB5_NOT_NOT)

LB1_NOT_NOT 3_NOT_NOT 1_NOT_NOT LB1_NOT_NOT
LB2_NOT_NOT 6_NOT_NOT 4_NOT_NOT LB2_NOT_NOT
LB3_NOT_NOT 8_NOT_NOT 9_NOT_NOT LB3_NOT_NOT
LB4_NOT_NOT 13_NOT_NOT 15_NOT_NOT LB4_NOT_NOT
LB5_NOT_NOT 21_NOT_NOT 23_NOT_NOT LB5_NOT_NOT

L1_NOT_NOT A_NOT_NOT 1_NOT_NOT 2.062E-12
L2_NOT_NOT 1_NOT_NOT 4_NOT_NOT 1.889E-12
L3_NOT_NOT 4_NOT_NOT 7_NOT_NOT 2.72E-12
L4_NOT_NOT CLK_NOT_NOT 13_NOT_NOT 2.057E-12
L5_NOT_NOT 13_NOT_NOT 16_NOT_NOT 1.029E-12
L6_NOT_NOT 16_NOT_NOT 17_NOT_NOT 1.241E-12
L7_NOT_NOT 16_NOT_NOT 12_NOT_NOT 1.973E-12
L8_NOT_NOT 10_NOT_NOT 12_NOT_NOT 1.003E-12
L9_NOT_NOT 10_NOT_NOT 8_NOT_NOT 7.524E-12
L10_NOT_NOT 8_NOT_NOT 20_NOT_NOT 1.234E-12
L11_NOT_NOT 18_NOT_NOT 21_NOT_NOT 2.607E-12
L12_NOT_NOT 21_NOT_NOT Q_NOT_NOT 2.062E-12

LP1_NOT_NOT 2_NOT_NOT 0 5.271E-13
LP2_NOT_NOT 5_NOT_NOT 0 5.237E-13
LP4_NOT_NOT 14_NOT_NOT 0 4.759E-13
LP6_NOT_NOT 11_NOT_NOT 0 5.021E-13
LP8_NOT_NOT 19_NOT_NOT 0 6.33E-13
LP9_NOT_NOT 22_NOT_NOT 0 4.749E-13

RB1_NOT_NOT 1_NOT_NOT 101_NOT_NOT RB1_NOT_NOT
LRB1_NOT_NOT 101_NOT_NOT 0 LRB1_NOT_NOT
RB2_NOT_NOT 4_NOT_NOT 104_NOT_NOT RB2_NOT_NOT
LRB2_NOT_NOT 104_NOT_NOT 5_NOT_NOT LRB2_NOT_NOT
RB3_NOT_NOT 7_NOT_NOT 107_NOT_NOT RB3_NOT_NOT
LRB3_NOT_NOT 107_NOT_NOT 8_NOT_NOT LRB3_NOT_NOT
RB4_NOT_NOT 13_NOT_NOT 113_NOT_NOT RB4_NOT_NOT
LRB4_NOT_NOT 113_NOT_NOT 0 LRB4_NOT_NOT
RB5_NOT_NOT 17_NOT_NOT 117_NOT_NOT RB5_NOT_NOT
LRB5_NOT_NOT 117_NOT_NOT 18_NOT_NOT LRB5_NOT_NOT
RB6_NOT_NOT 10_NOT_NOT 110_NOT_NOT RB6_NOT_NOT
LRB6_NOT_NOT 110_NOT_NOT 0 LRB6_NOT_NOT
RB7_NOT_NOT 20_NOT_NOT 120_NOT_NOT RB7_NOT_NOT
LRB7_NOT_NOT 120_NOT_NOT 18_NOT_NOT LRB7_NOT_NOT
RB8_NOT_NOT 18_NOT_NOT 118_NOT_NOT RB8_NOT_NOT
LRB8_NOT_NOT 118_NOT_NOT 0 LRB8_NOT_NOT
RB9_NOT_NOT 21_NOT_NOT 121_NOT_NOT RB9_NOT_NOT
LRB9_NOT_NOT 121_NOT_NOT 0 LRB9_NOT_NOT
LRD_NOT_NOT 12_NOT_NOT 112_NOT_NOT LRD_NOT_NOT
RD_NOT_NOT 112_NOT_NOT 0 RD_NOT_NOT




*JTL_NOT

LC_JTL_NOT_1 CLKD A_JTL_NOT 0
LC_JTL_NOT_2 CLK Q_JTL_NOT 0

.MODEL JJMIT_JTL_NOT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.PARAM PHI0_JTL_NOT = 2.0678E-15
.PARAM B0_JTL_NOT = 1
.PARAM IC0_JTL_NOT = 1.0000E-04
.PARAM ICRS_JTL_NOT = 6.8599E-04
.PARAM B0RS_JTL_NOT = 6.8599
.PARAM RSHEET_JTL_NOT = 2
.PARAM LSHEET_JTL_NOT = 1.1300E-12
.PARAM LP_JTL_NOT = 2.0000E-13
.PARAM IC_JTL_NOT = 2.5000
.PARAM LPTL_JTL_NOT = 2.0000E-12
.PARAM LB_JTL_NOT = 2.0000E-12
.PARAM BIASCOEF_JTL_NOT = 0.7000
.PARAM B1_JTL_NOT = 2.5000
.PARAM B2_JTL_NOT = 2.5000
.PARAM IB1_JTL_NOT = 3.5000E-04
.PARAM LB1_JTL_NOT = 2.0000E-12
.PARAM L1_JTL_NOT = 2.0678E-12
.PARAM L2_JTL_NOT = 2.0678E-12
.PARAM L3_JTL_NOT = 2.0678E-12
.PARAM L4_JTL_NOT = 2.0678E-12
.PARAM RB1_JTL_NOT = 2.7440
.PARAM RB2_JTL_NOT = 2.7440
.PARAM LRB1_JTL_NOT = 1.7503E-12
.PARAM LRB2_JTL_NOT = 1.7503E-12
.PARAM LP1_JTL_NOT = 2.0000E-13
.PARAM LP2_JTL_NOT = 2.0000E-13

B1_JTL_NOT 1_JTL_NOT 2_JTL_NOT JJMIT_JTL_NOT AREA=B1_JTL_NOT
B2_JTL_NOT 6_JTL_NOT 7_JTL_NOT JJMIT_JTL_NOT AREA=B2_JTL_NOT
IB1_JTL_NOT 0 5_JTL_NOT PWL(0 0 5P IB1_JTL_NOT)
L1_JTL_NOT A_JTL_NOT 1_JTL_NOT 2.082E-12
L2_JTL_NOT 1_JTL_NOT 4_JTL_NOT 2.06E-12
L3_JTL_NOT 4_JTL_NOT 6_JTL_NOT 2.067E-12
L4_JTL_NOT 6_JTL_NOT Q_JTL_NOT 2.075E-12
LP1_JTL_NOT 2_JTL_NOT 0 4.998E-13
LP2_JTL_NOT 7_JTL_NOT 0 5.011E-13
LB1_JTL_NOT 5_JTL_NOT 4_JTL_NOT LB1_JTL_NOT
RB1_JTL_NOT 1_JTL_NOT 3_JTL_NOT RB1_JTL_NOT
RB2_JTL_NOT 6_JTL_NOT 8_JTL_NOT RB2_JTL_NOT
LRB1_JTL_NOT 3_JTL_NOT 0 LRB1_JTL_NOT
LRB2_JTL_NOT 8_JTL_NOT 0 LRB2_JTL_NOT


*OR_NOT

LC_OR_NOT_1 BNNN A_OR_NOT 0
LC_OR_NOT_2 CNNN B_OR_NOT 0
LC_OR_NOT_3 CLKD Q_OR_NOT 0

* .SUBCKT DSFQ_OR_NOT A_OR_NOT B_OR_NOT Q_OR_NOT
.MODEL JJMIT_OR_NOT JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
*CONFLUENCE BUFFER A
.PARAM L1_OR_NOT = 2E-12
.PARAM B1_OR_NOT = 1.37211310E+00
.PARAM B3_OR_NOT = 2.77209629E+00
.PARAM B4_OR_NOT = 3.78734058E-01

* AND GATE LOOP
.PARAM L4_OR_NOT = 1.22182342E-12
.PARAM B7_OR_NOT = 1.19265113E+00
.PARAM B9_OR_NOT = 5.40924075E-01
.PARAM L7_OR_NOT = 1.62539785E-13
.PARAM R1_OR_NOT = 1.09745275E+01
.PARAM R2_OR_NOT = 5.58089917E-01
.PARAM L5_OR_NOT = 5.61756493E-13

* OUTPUT STAGE
.PARAM B8_OR_NOT = 7.09413113E-01
.PARAM I1_OR_NOT = 3.23631555E-04
.PARAM L3_OR_NOT = 2E-12
.PARAM L6_OR_NOT = 3.06315548E-12

*CONFLUENCE BUFFER B
.PARAM L2_OR_NOT = L1_OR_NOT
.PARAM B2_OR_NOT = B1_OR_NOT
.PARAM B5_OR_NOT = B3_OR_NOT
.PARAM B6_OR_NOT = B4_OR_NOT

*PARASITICS
.PARAM LP1_OR_NOT = 0.2E-12
.PARAM LP2_OR_NOT = 0.2E-12
.PARAM LP3_OR_NOT = 0.2E-12
.PARAM LP4_OR_NOT = 0.2E-12

* BACK ANNOTATED .CIR FILE FROM KICAD
B1_OR_NOT 3_OR_NOT 1_OR_NOT JJMIT_OR_NOT AREA=B1_OR_NOT
B2_OR_NOT 4_OR_NOT 2_OR_NOT JJMIT_OR_NOT AREA=B2_OR_NOT
B3_OR_NOT 3_OR_NOT 10_OR_NOT JJMIT_OR_NOT AREA=B3_OR_NOT
B4_OR_NOT 5_OR_NOT 3_OR_NOT JJMIT_OR_NOT AREA=B4_OR_NOT
B5_OR_NOT 4_OR_NOT 10_OR_NOT JJMIT_OR_NOT AREA=B5_OR_NOT
B6_OR_NOT 6_OR_NOT 4_OR_NOT JJMIT_OR_NOT AREA=B6_OR_NOT
B7_OR_NOT 24_OR_NOT 20_OR_NOT JJMIT_OR_NOT AREA=B7_OR_NOT
B8_OR_NOT 30_OR_NOT 31_OR_NOT JJMIT_OR_NOT AREA=B8_OR_NOT
B9_OR_NOT 24_OR_NOT 23_OR_NOT JJMIT_OR_NOT AREA=B9_OR_NOT
I1_OR_NOT 0 10_OR_NOT PWL(0 0 5P I1_OR_NOT)
L1_OR_NOT A_OR_NOT 1_OR_NOT L1_OR_NOT
L2_OR_NOT B_OR_NOT 2_OR_NOT L2_OR_NOT
L3_OR_NOT 10_OR_NOT 30_OR_NOT L3_OR_NOT
L4_OR_NOT 30_OR_NOT 20_OR_NOT L4_OR_NOT
L5_OR_NOT 21_OR_NOT 24_OR_NOT L5_OR_NOT
L6_OR_NOT 30_OR_NOT Q_OR_NOT L6_OR_NOT
L7_OR_NOT 22_OR_NOT 23_OR_NOT L7_OR_NOT
LP1_OR_NOT 5_OR_NOT 0 LP1_OR_NOT
LP2_OR_NOT 6_OR_NOT 0 LP2_OR_NOT
LP3_OR_NOT 24_OR_NOT 0 LP3_OR_NOT
LP4_OR_NOT 31_OR_NOT 0 LP4_OR_NOT
R1_OR_NOT 21_OR_NOT 20_OR_NOT R1_OR_NOT
R2_OR_NOT 22_OR_NOT 20_OR_NOT R2_OR_NOT


*** SPLIT CELLS********************************************************************************************************************************

LC_SPLIT1_1 A A_SPLIT1 0
LC_SPLIT1_2 A1 Q0_SPLIT1 0
LC_SPLIT1_3 A2 Q1_SPLIT1 0
.MODEL JJMIT_SPLIT1 JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.PARAM PHI0_SPLIT1 = 2.0678E-15
.PARAM B0_SPLIT1 = 1
.PARAM IC0_SPLIT1 = 1.0000E-04
.PARAM ICRS_SPLIT1 = 6.8599E-04
.PARAM B0RS_SPLIT1 = 6.8599
.PARAM RSHEET_SPLIT1 = 2
.PARAM LSHEET_SPLIT1 = 1.1300E-12
.PARAM LP_SPLIT1 = 2.0000E-13
.PARAM IC_SPLIT1 = 2.5000
.PARAM LPTL_SPLIT1 = 2.0000E-12
.PARAM LB_SPLIT1 = 2.0000E-12
.PARAM BIASCOEF_SPLIT1 = 0.7000
.PARAM RD_SPLIT1 = 1.3600
.PARAM B1_SPLIT1 = 2.5000
.PARAM B2_SPLIT1 = 3
.PARAM B3_SPLIT1 = 2.5000
.PARAM B4_SPLIT1 = 2.5000
.PARAM IB1_SPLIT1 = 1.7500E-04
.PARAM IB2_SPLIT1 = 2.8000E-04
.PARAM IB3_SPLIT1 = 1.7500E-04
.PARAM IB4_SPLIT1 = 1.7500E-04
.PARAM L1_SPLIT1 = 2.0000E-12
.PARAM L2_SPLIT1 = 4.1357E-12
.PARAM L3_SPLIT1 = 1.7232E-12
.PARAM L4_SPLIT1 = 1.7232E-12
.PARAM L5_SPLIT1 = 2.0000E-12
.PARAM L6_SPLIT1 = 1.7232E-12
.PARAM L7_SPLIT1 = 2.0000E-12
.PARAM RB1_SPLIT1 = 2.7440
.PARAM RB2_SPLIT1 = 2.2866
.PARAM RB3_SPLIT1 = 2.7440
.PARAM RB4_SPLIT1 = 2.7440
.PARAM LRB1_SPLIT1 = 1.5503E-12
.PARAM LRB2_SPLIT1 = 1.2919E-12
.PARAM LRB3_SPLIT1 = 1.5503E-12
.PARAM LRB4_SPLIT1 = 1.5503E-12

IB1_SPLIT1 0 3_SPLIT1 PWL(0 0 5P IB1_SPLIT1)
IB2_SPLIT1 0 6_SPLIT1 PWL(0 0 5P IB2_SPLIT1)
IB3_SPLIT1 0 10_SPLIT1 PWL(0 0 5P IB3_SPLIT1)
IB4_SPLIT1 0 13_SPLIT1 PWL(0 0 5P IB4_SPLIT1)
LB1_SPLIT1 3_SPLIT1 1_SPLIT1 9.175E-13
LB2_SPLIT1 6_SPLIT1 4_SPLIT1 7.666E-13
LB3_SPLIT1 10_SPLIT1 8_SPLIT1 1.928E-12
LB4_SPLIT1 13_SPLIT1 11_SPLIT1 8.786E-13

B1_SPLIT1 1_SPLIT1 2_SPLIT1 JJMIT_SPLIT1 AREA=B1_SPLIT1
B2_SPLIT1 4_SPLIT1 5_SPLIT1 JJMIT_SPLIT1 AREA=B2_SPLIT1
B3_SPLIT1 8_SPLIT1 9_SPLIT1 JJMIT_SPLIT1 AREA=B3_SPLIT1
B4_SPLIT1 11_SPLIT1 12_SPLIT1 JJMIT_SPLIT1 AREA=B4_SPLIT1
L1_SPLIT1 A_SPLIT1 1_SPLIT1 2.063E-12
L2_SPLIT1 1_SPLIT1 4_SPLIT1 3.637E-12
L3_SPLIT1 4_SPLIT1 7_SPLIT1 1.278E-12
L4_SPLIT1 7_SPLIT1 8_SPLIT1 1.305E-12
L5_SPLIT1 8_SPLIT1 Q0_SPLIT1 2.05E-12
L6_SPLIT1 7_SPLIT1 11_SPLIT1 1.315E-12
L7_SPLIT1 11_SPLIT1 Q1_SPLIT1 2.06E-12

LP1_SPLIT1 2_SPLIT1 0 4.676E-13
LP2_SPLIT1 5_SPLIT1 0 4.498E-13
LP3_SPLIT1 9_SPLIT1 0 5.183E-13
LP4_SPLIT1 12_SPLIT1 0 4.639E-13
RB1_SPLIT1 1_SPLIT1 101_SPLIT1 RB1_SPLIT1
LRB1_SPLIT1 101_SPLIT1 0 LRB1_SPLIT1
RB2_SPLIT1 4_SPLIT1 104_SPLIT1 RB2_SPLIT1
LRB2_SPLIT1 104_SPLIT1 0 LRB2_SPLIT1
RB3_SPLIT1 8_SPLIT1 108_SPLIT1 RB3_SPLIT1
LRB3_SPLIT1 108_SPLIT1 0 LRB3_SPLIT1
RB4_SPLIT1 11_SPLIT1 111_SPLIT1 RB4_SPLIT1
LRB4_SPLIT1 111_SPLIT1 0 LRB4_SPLIT1



*SPLIT2



LC_SPLIT2_1 B A_SPLIT2 0
LC_SPLIT2_2 B1 Q0_SPLIT2 0
LC_SPLIT2_3 B2 Q1_SPLIT2 0
.MODEL JJMIT_SPLIT2 JJ(RTYPE=1, VG=2.8MV, CAP=0.07PF, R0=160, RN=16, ICRIT=0.1MA)
.PARAM PHI0_SPLIT2 = 2.0678E-15
.PARAM B0_SPLIT2 = 1
.PARAM IC0_SPLIT2 = 1.0000E-04
.PARAM ICRS_SPLIT2 = 6.8599E-04
.PARAM B0RS_SPLIT2 = 6.8599
.PARAM RSHEET_SPLIT2 = 2
.PARAM LSHEET_SPLIT2 = 1.1300E-12
.PARAM LP_SPLIT2 = 2.0000E-13
.PARAM IC_SPLIT2 = 2.5000
.PARAM LPTL_SPLIT2 = 2.0000E-12
.PARAM LB_SPLIT2 = 2.0000E-12
.PARAM BIASCOEF_SPLIT2 = 0.7000
.PARAM RD_SPLIT2 = 1.3600
.PARAM B1_SPLIT2 = 2.5000
.PARAM B2_SPLIT2 = 3
.PARAM B3_SPLIT2 = 2.5000
.PARAM B4_SPLIT2 = 2.5000
.PARAM IB1_SPLIT2 = 1.7500E-04
.PARAM IB2_SPLIT2 = 2.8000E-04
.PARAM IB3_SPLIT2 = 1.7500E-04
.PARAM IB4_SPLIT2 = 1.7500E-04
.PARAM L1_SPLIT2 = 2.0000E-12
.PARAM L2_SPLIT2 = 4.1357E-12
.PARAM L3_SPLIT2 = 1.7232E-12
.PARAM L4_SPLIT2 = 1.7232E-12
.PARAM L5_SPLIT2 = 2.0000E-12
.PARAM L6_SPLIT2 = 1.7232E-12
.PARAM L7_SPLIT2 = 2.0000E-12
.PARAM RB1_SPLIT2 = 2.7440
.PARAM RB2_SPLIT2 = 2.2866
.PARAM RB3_SPLIT2 = 2.7440
.PARAM RB4_SPLIT2 = 2.7440
.PARAM LRB1_SPLIT2 = 1.5503E-12
.PARAM LRB2_SPLIT2 = 1.2919E-12
.PARAM LRB3_SPLIT2 = 1.5503E-12
.PARAM LRB4_SPLIT2 = 1.5503E-12

IB1_SPLIT2 0 3_SPLIT2 PWL(0 0 5P IB1_SPLIT2)
IB2_SPLIT2 0 6_SPLIT2 PWL(0 0 5P IB2_SPLIT2)
IB3_SPLIT2 0 10_SPLIT2 PWL(0 0 5P IB3_SPLIT2)
IB4_SPLIT2 0 13_SPLIT2 PWL(0 0 5P IB4_SPLIT2)
LB1_SPLIT2 3_SPLIT2 1_SPLIT2 9.175E-13
LB2_SPLIT2 6_SPLIT2 4_SPLIT2 7.666E-13
LB3_SPLIT2 10_SPLIT2 8_SPLIT2 1.928E-12
LB4_SPLIT2 13_SPLIT2 11_SPLIT2 8.786E-13

B1_SPLIT2 1_SPLIT2 2_SPLIT2 JJMIT_SPLIT2 AREA=B1_SPLIT2
B2_SPLIT2 4_SPLIT2 5_SPLIT2 JJMIT_SPLIT2 AREA=B2_SPLIT2
B3_SPLIT2 8_SPLIT2 9_SPLIT2 JJMIT_SPLIT2 AREA=B3_SPLIT2
B4_SPLIT2 11_SPLIT2 12_SPLIT2 JJMIT_SPLIT2 AREA=B4_SPLIT2
L1_SPLIT2 A_SPLIT2 1_SPLIT2 2.063E-12
L2_SPLIT2 1_SPLIT2 4_SPLIT2 3.637E-12
L3_SPLIT2 4_SPLIT2 7_SPLIT2 1.278E-12
L4_SPLIT2 7_SPLIT2 8_SPLIT2 1.305E-12
L5_SPLIT2 8_SPLIT2 Q0_SPLIT2 2.05E-12
L6_SPLIT2 7_SPLIT2 11_SPLIT2 1.315E-12
L7_SPLIT2 11_SPLIT2 Q1_SPLIT2 2.06E-12

LP1_SPLIT2 2_SPLIT2 0 4.676E-13
LP2_SPLIT2 5_SPLIT2 0 4.498E-13
LP3_SPLIT2 9_SPLIT2 0 5.183E-13
LP4_SPLIT2 12_SPLIT2 0 4.639E-13
RB1_SPLIT2 1_SPLIT2 101_SPLIT2 RB1_SPLIT2
LRB1_SPLIT2 101_SPLIT2 0 LRB1_SPLIT2
RB2_SPLIT2 4_SPLIT2 104_SPLIT2 RB2_SPLIT2
LRB2_SPLIT2 104_SPLIT2 0 LRB2_SPLIT2
RB3_SPLIT2 8_SPLIT2 108_SPLIT2 RB3_SPLIT2
LRB3_SPLIT2 108_SPLIT2 0 LRB3_SPLIT2
RB4_SPLIT2 11_SPLIT2 111_SPLIT2 RB4_SPLIT2
LRB4_SPLIT2 111_SPLIT2 0 LRB4_SPLIT2

* .ENDS

.ends