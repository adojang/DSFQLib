.title KiCad schematic
LRB5 /32 GND Inductor
LP1 /31 GND Inductor
LRB4 Net-_LRB4-Pad1_ /30 Inductor
RB4 /22 Net-_LRB4-Pad1_ Resistor
B5 /31 /30 jjmit
RB3 /12 Net-_LRB3-Pad1_ Resistor
LRB3 Net-_LRB3-Pad1_ /30 Inductor
L3 /30 Q Inductor
RB5 /30 /32 Resistor
I1 GND /30 pwl(0 0 5p REF)
L2 B /20 Inductor
B1 /30 /10 jjmit
R1 /10 /30 Resistor
R3 /12 /10 Resistor
LRB1 /11 /30 Inductor
RB1 /10 /11 Resistor
B3 /30 /12 jjmit
R2 /20 /30 Resistor
B2 /30 /20 jjmit
B4 /30 /22 jjmit
RB2 /20 /21 Resistor
LRB2 /21 /30 Inductor
R4 /22 /20 Resistor
L1 A /10 Inductor
.end
