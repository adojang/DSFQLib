.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_SFQDC_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include AW_mitll_DSFQ_AND.cir

.tran 0.015p 250p 0
.param cval= 600u

*15ps skew with 2e-12 input.
I_A0 0 xa pwl(0 0 100p 0 103p cval 105p 0)
* I_A1 0 xc pwl(0 0 100p 0 103p cval 105p 0 200p 0 203p 0 205p 0) 
* I_B1 0 xd pwl(0 0 100p 0 103p cval 105p 0 213p cval 216p 0 218p 0)

XDCSFQA LSmitll_DCSFQ xa xa1 

* XDCSFQC LSmitll_DCSFQ xc xc1 
* XDCSFQD LSmitll_DCSFQ xd xd1


XJTLA LSMITLL_JTL xa1 A

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)


L1      A       B       7p
RH      B       Ba      4
LHp     Ba      Q       0.5p
BS      B       Q       jjmit area=0.84
BD      C       Q       jjmit area=0.6
RD      B       Bb      0.68
LDp     Bb      C       0.5p

.print p(A) i(L1) i(BS) p(Q) 




*Print Full Phase for Appendix

XLOAD LSMITLL_JTL q qq

Rsink qq 0 2
