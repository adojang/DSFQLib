.title KiCad schematic
L6 /12 /13 Inductor
L7 /13 /16 Inductor
B6 /12 /4 jjmit
B9 /15 /17 jjmit
LP5 /15 GND Inductor
LP4 /14 GND Inductor
B8 /14 /13 jjmit
I3 GND /16 pwl(0 0 5p REF)
L8 /16 /17 Inductor
L9 /17 Q Inductor
B7 /8 /12 jjmit
LP3 /8 GND Inductor
L10 /102 /104 Inductor
L5 A /101 Inductor
B10 /102 /101 jjmit
B2 /6 /5 jjmit
B11 /103 /102 jjmit
LP6 /103 GND Inductor
L1 CLK /55 Inductor
L11 /104 /105 Inductor
I4 unconnected-_I4-Pad1_ /104 pwl(0 0 5p REF)
B1 /5 /55 jjmit
B5 /4 /44 jjmit
B12 /106 /105 jjmit
L12 /105 /44 Inductor
LP7 /106 GND Inductor
B4 /12 /11 jjmit
L4 /10 /11 Inductor
I2 GND /4 pwl(0 0 5p REF)
L3 /9 /10 Inductor
I1 GND /9 pwl(0 0 5p REF)
L2 /5 /9 Inductor
LP2 /7 GND Inductor
B3 /7 /10 jjmit
LP1 /6 GND Inductor
.end
