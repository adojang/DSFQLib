.subckt DSFQ_INV A CLK Q

.param b3  =	         0.975397461
.param b4  =	         1.97590602
.param b5  =	         6.82124243e-01
.param b6  =	         2.77586674e-01
.param b7 =	 	       5.35250160e-01
.param b8 =	 	       5.98173295e-01
.param b9 =	 	       1.22329715e+00
.param i1 =	 	       1.18063229e-04
.param i2 =	 	       6.31851665e-05
.param i3 =	 	       1.04993869e-04
.param l10  =    1.78304590e-12
.param l2  =     1.76930775e-12
.param l3  =     1.77358790e-12
.param l4  =     1.45997109e-12
.param l5  =     1.77468740e-12
.param l6  =     2.48124061e-12
.param l7  =     1.46863740e-12
.param l8  =     1.46042354e-12
.param l9  =     1.46832533e-12
.param 	lp1  	= 0.2p
.param 	lp2  	= 0.2p
.param 	lp3  	= 0.2p
.param 	lp4  	= 0.2p
.param 	lp5  	= 0.2p


* Back Annotated .cir file from KiCad
b3   	12   	4   	 jjmit area=b3
b4   	12   	11   	 jjmit area=b4
b5   	6   	5   	 jjmit area=b5
b6   	7   	10   	 jjmit area=b6
b7   	14   	13   	 jjmit area=b7
b8   	15   	17   	 jjmit area=b8
b9   	8   	12   	 jjmit area=b9
i1   	0   	9   	pwl(0   	0   	5p   	i1)
i2   	0   	16   	pwl(0   	0   	5p   	i2)
i3   	0   	4   	pwl(0   	0   	5p   	i3)
l10   	17   	Q   	 l10
l2   	A   	4   	 l2
l3   	CLK   	5   	 l3
l4   	5   	9   	 l4
l5   	9   	10   	 l5
l6   	10   	11   	 l6
l7   	12   	13   	 l7
l8   	13   	16   	 l8
l9   	16   	17   	 l9
lp1   	6   	0   	 lp1
lp2   	7   	0   	 lp2
lp3   	14   	0   	 lp3
lp4   	15   	0   	 lp4
lp5   	8   	0   	 lp5
.ends