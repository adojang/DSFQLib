1.6874e-10      0     0     0     1        0
2.6822e-10      1     0     0     1        0
3.6874e-10      1     0     1     1        0
4.6874e-10      2     1     1     1        0 # THIS INDEX
5.6826e-10      2     1     1     2        0
6.6826e-10      2     1     2     2        0
7.6827e-10      2     1     3     3        0
8.687e-10       3     1     3     3        0
1.06874e-09     3     2     3     3        0
1.16828e-09     4     3     3     3        0
1.26827e-09     4     4     3     3        0
1.36874e-09     4     4     4     4        0


if 4 == 4 then set new == 0
if 5 > 4 set new == 1

if a == b set new = 0
if a != b set new = 1

Desired OUTPUT:

00010
10000
00101
11000