.subckt DSFQ_MUX D0 D1 S QQ

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)

.param B2 = 0.8
.param Q2 = 0.8
.param A2 = 0.8
.param A1 = 3.35

B_x2   B2   	0   	 jjmit area=B2
B_xQ2  	Q2x   	0   	 jjmit area=Q2
B_xA2  	A2   	0   	 jjmit area=A2
B_xA1   A1   	0   	 jjmit area=A1

XSPLITA LSMITLL_SPLITm D0 A1x CLKx
XSPLITB LSMITLL_SPLITm D1 B1x B1x
XSPLITS LSMITLL_SPLITm S S1x B2x

XCJTLA1 LSMITLL_JTLm A1x A1
XCJTLA2 LSMITLL_JTLm A2x A2
XCJTLCLK LSMITLL_JTLm CLKx CLK
XCJTLS1 LSMITLL_JTLm S1x S1
XCJTLB1 LSMITLL_JTLm B1x B1
XCJTLB2 LSMITLL_JTLm B2x B2

XQ1 LSMITLL_JTLm Q1x Q1
XQ2 LSMITLL_JTLm Q2x Q2


XAND1   DSFQ_ANDm   A1 A2 Q1x
XAND2   DSFQ_ANDm   B1 B2 Q2x
XNOT    DSFQ_NOTm S1 CLK CLK A2x
XOR     DSFQ_ORm    Q1 Q2 QQ




* Back-annotated simulation file written by InductEx v.6.0.4 on 1-4-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 9 March 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

* The cell is not designed to be connected directly to passive transmission lines

*$Ports a q0 q1
.subckt LSmitll_SPLITm a q0 q1
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7
.param RD=1.36

.param B1=2.5
.param B2=3.0
.param B3=2.5
.param B4=2.5

.param IB1=175u
.param IB2=280u
.param IB3=175u
.param IB4=175u

.param L1=Lptl
.param L2=Phi0/(2*B1*Ic0)
.param L3=(Phi0/(2*B2*Ic0))/2
.param L4=L3
.param L5=Lptl
.param L6=L3
.param L7=Lptl

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 10 pwl(0 0 5p IB3)
IB4 0 13 pwl(0 0 5p IB4)
LB1 3 1 9.175E-13
LB2 6 4 7.666E-13
LB3 10 8 1.928E-12
LB4 13 11 8.786E-13

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 8 9 jjmit area=B3
B4 11 12 jjmit area=B4
L1 a 1 2.063E-12
L2 1 4 3.637E-12
L3 4 7 1.278E-12
L4 7 8 1.305E-12
L5 8 q0 2.05E-12
L6 7 11 1.315E-12
L7 11 q1 2.06E-12

LP1 2 0 4.676E-13
LP2 5 0 4.498E-13
LP3 9 0 5.183E-13
LP4 12 0 4.639E-13
RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 0 LRB2
RB3 8 108 RB3
LRB3 108 0 LRB3
RB4 11 111 RB4
LRB4 111 0 LRB4
.ends



* Back-annotated simulation file written by InductEx v.6.0.4 on 10-3-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 12 January 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

* The cell is not designed to be connected directly to passive transmission lines

*$Ports 			a q
.subckt LSMITLL_JTLm a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=IC
.param IB1=(B1+B2)*Ic0*BiasCoef
.param LB1=LB
.param L1=Phi0/(4*B1*Ic0)
.param L2=Phi0/(4*B1*Ic0)
.param L3=Phi0/(4*B1*Ic0)
.param L4=Phi0/(4*B2*Ic0)
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP

B1 1 2 jjmit area=B1
B2 6 7 jjmit area=B2
IB1 0 5 pwl(0 0 5p IB1)
L1 a 1 2.082E-12
L2 1 4 2.06E-12
L3 4 6 2.067E-12
L4 6 q 2.075E-12
LP1 2 0 4.998E-13
LP2 7 0 5.011E-13
LB1 5 4 LB1
RB1 1 3 RB1
RB2 6 8 RB2
LRB1 3 0 LRB1
LRB2 8 0 LRB2
.ends



.subckt DSFQ_ANDm A B Q
.param b1  	=	 1.39878486e+00
.param bd1  =	 1.38855937e+00
.param l1  	=	 2e-12
.param rd1  =	 6.00718616e-01
.param i1  	=	 1.54457273e-05
.param b3  	=	 1.51517089e+00
.param l3  	=	 2e-12
.param rh1  =	 4.76237371e+00

*Parasitics and Matching
.param 	ldp1  	= 1e-12
.param 	b2  	= b1
.param 	bd2  	= bd1
.param 	l2  	= l1
.param 	ldp2  	= ldp1
.param 	rd2  	= rd1
.param 	lp1  	= 0.2e-12
.param 	lhp1  	= 1e-12
.param 	lhp2  	= lhp1
.param 	rh2  	= rh1

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

* Back Annotated .cir file from KiCad
b1   	30   	10   	 jjmit area=b1
b2   	30   	20   	 jjmit area=b2
b3   	31   	30   	 jjmit area=b3
bd1   	30   	12   	 jjmit area=bd1
bd2   	30   	22   	 jjmit area=bd2
i1   	0   	30   	pwl(0   	0   	5p   	i1)
l1   	a   	10   	 l1
l2   	b   	20   	 l2
l3   	30   	q   	 l3
ldp1   	11   	12   	 ldp1
ldp2   	21   	22   	 ldp2
lhp1   	13   	30   	 lhp1
lhp2   	23   	30   	 lhp2
lp1   	31   	0   	 lp1
rd1   	11   	10   	 rd1
rd2   	21   	20   	 rd2
rh1   	13   	10   	 rh1
rh2   	23   	20   	 rh2
.ends

.subckt DSFQ_NOTm A B C Q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
*A is inverting input.
*B and C are inputs for the OR gate.
*Q is output.

XDSFQ_OR DSFQ_ORi B C CLKD
XJTLCLK LSMITLL_JTLi CLKD CLK
XNOTLS LSMITLL_NOTi A CLK Q



.subckt DSFQ_ORi a b q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
*Confluence Buffer A
.param l1  	=	 	    2e-12
.param b1  	=	 	    1.37211310e+00
.param b3  	=	 	    2.77209629e+00
.param b4  	=	 	    3.78734058e-01

* AND GATE LOOP
.param l4  	=	 	    1.22182342e-12
.param b7  	=	 	    1.19265113e+00
.param b9  	=	 	    5.40924075e-01
.param l7  	=	 	    1.62539785e-13
.param r1  	=	 	    1.09745275e+01
.param r2  	=	 	    5.58089917e-01
.param l5  	=	 	    5.61756493e-13

* Output Stage
.param b8  	=	 	    7.09413113e-01
.param i1  	=	 	    3.23631555e-04
.param l3  	=	 	   2e-12
.param l6  	=	 	    3.06315548e-12

*Confluence Buffer B
.param 	l2  	= L1
.param 	b2  	= B1
.param 	b5  	= B3
.param 	b6  	= B4

*Parasitics
.param 	lp1  	= 0.2e-12
.param 	lp2  	= 0.2e-12
.param 	lp3  	= 0.2e-12
.param 	lp4  	= 0.2e-12

* Back Annotated .cir file from KiCad
b1   	3   	1   	 jjmit area=b1
b2   	4   	2   	 jjmit area=b2
b3   	3   	10   	 jjmit area=b3
b4   	5   	3   	 jjmit area=b4
b5   	4   	10   	 jjmit area=b5
b6   	6   	4   	 jjmit area=b6
b7   	24   	20   	 jjmit area=b7
b8   	30   	31   	 jjmit area=b8
b9   	24   	23   	 jjmit area=b9
i1   	0   	10   	pwl(0   	0   	5p      i1)
l1   	a   	1   	 l1
l2   	b   	2   	 l2
l3   	10   	30   	 l3
l4   	30   	20   	 l4
l5   	21   	24   	 l5
l6   	30   	q   	 l6
l7   	22   	23   	 l7
lp1   	5   	0   	 lp1
lp2   	6   	0   	 lp2
lp3   	24   	0   	 lp3
lp4   	31   	0   	 lp4
r1   	21   	20   	 r1
r2   	22   	20   	 r2
.ends



.subckt DSFQ_ORm a b q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
*Confluence Buffer A
.param l1  	=	 	    2e-12
.param b1  	=	 	    1.37211310e+00
.param b3  	=	 	    2.77209629e+00
.param b4  	=	 	    3.78734058e-01

* AND GATE LOOP
.param l4  	=	 	    1.22182342e-12
.param b7  	=	 	    1.19265113e+00
.param b9  	=	 	    5.40924075e-01
.param l7  	=	 	    1.62539785e-13
.param r1  	=	 	    1.09745275e+01
.param r2  	=	 	    5.58089917e-01
.param l5  	=	 	    5.61756493e-13

* Output Stage
.param b8  	=	 	    7.09413113e-01
.param i1  	=	 	    3.23631555e-04
.param l3  	=	 	    2e-12
.param l6  	=	 	    3.06315548e-12

*Confluence Buffer B
.param 	l2  	= L1
.param 	b2  	= B1
.param 	b5  	= B3
.param 	b6  	= B4

*Parasitics
.param 	lp1  	= 0.2e-12
.param 	lp2  	= 0.2e-12
.param 	lp3  	= 0.2e-12
.param 	lp4  	= 0.2e-12

* Back Annotated .cir file from KiCad
b1   	3   	1   	 jjmit area=b1
b2   	4   	2   	 jjmit area=b2
b3   	3   	10   	 jjmit area=b3
b4   	5   	3   	 jjmit area=b4
b5   	4   	10   	 jjmit area=b5
b6   	6   	4   	 jjmit area=b6
b7   	24   	20   	 jjmit area=b7
b8   	30   	31   	 jjmit area=b8
b9   	24   	23   	 jjmit area=b9
i1   	0   	10   	pwl(0   	0   	5p      i1)
l1   	a   	1   	 l1
l2   	b   	2   	 l2
l3   	10   	30   	 l3
l4   	30   	20   	 l4
l5   	21   	24   	 l5
l6   	30   	q   	 l6
l7   	22   	23   	 l7
lp1   	5   	0   	 lp1
lp2   	6   	0   	 lp2
lp3   	24   	0   	 lp3
lp4   	31   	0   	 lp4
r1   	21   	20   	 r1
r2   	22   	20   	 r2
.ends



* Back-annotated simulation file written by InductEx v.6.0.4 on 8-4-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 3 June 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

* The cell is not designed to be connected directly to passive transmission lines

*$Ports  a clk q
.subckt LSMITLL_NOTi a clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=2.57
.param B3=1.07
.param B4=IC
.param B5=1.34
.param B6=3.03
.param B7=1.38
.param B8=0.8
.param B9=IC

.param IB1=BiasCoef*Ic0*B1
.param IB2=87u
.param IB3=257u
.param IB4=BiasCoef*Ic0*B4
.param IB5=BiasCoef*Ic0*B9

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9

.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet

.param RD=4
.param LRD=2p

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 7 8 jjmit area=B3
B4 13 14 jjmit area=B4
B5 17 18 jjmit area=B5
B6 10 11 jjmit area=B6
B7 20 18 jjmit area=B7
B8 18 19 jjmit area=B8
B9 21 22 jjmit area=B9

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 9 pwl(0 0 5p IB3)
IB4 0 15 pwl(0 0 5p IB4)
IB5 0 23 pwl(0 0 5p IB5)

LB1 3 1 LB1
LB2 6 4 LB2
LB3 8 9 LB3
LB4 13 15 LB4
LB5 21 23 LB5

L1 a 1 2.062E-12
L2 1 4 1.889E-12
L3 4 7 2.72E-12
L4 clk 13 2.057E-12
L5 13 16 1.029E-12
L6 16 17 1.241E-12
L7 16 12 1.973E-12
L8 10 12 1.003E-12
L9 10 8 7.524E-12
L10 8 20 1.234E-12
L11 18 21 2.607E-12
L12 21 q 2.062E-12

LP1 2 0 5.271E-13
LP2 5 0 5.237E-13
LP4 14 0 4.759E-13
LP6 11 0 5.021E-13
LP8 19 0 6.33E-13
LP9 22 0 4.749E-13

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 5 LRB2
RB3 7 107 RB3
LRB3 107 8 LRB3
RB4 13 113 RB4
LRB4 113 0 LRB4
RB5 17 117 RB5
LRB5 117 18 LRB5
RB6 10 110 RB6
LRB6 110 0 LRB6
RB7 20 120 RB7
LRB7 120 18 LRB7
RB8 18 118 RB8
LRB8 118 0 LRB8
RB9 21 121 RB9
LRB9 121 0 LRB9
LRD 12 112 LRD
RD 112 0 RD
.ends

* Back-annotated simulation file written by InductEx v.6.0.4 on 10-3-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 12 January 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

* The cell is not designed to be connected directly to passive transmission lines

*$Ports 			a q
.subckt LSMITLL_JTLi a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=IC
.param IB1=(B1+B2)*Ic0*BiasCoef
.param LB1=LB
.param L1=Phi0/(4*B1*Ic0)
.param L2=Phi0/(4*B1*Ic0)
.param L3=Phi0/(4*B1*Ic0)
.param L4=Phi0/(4*B2*Ic0)
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP

B1 1 2 jjmit area=B1
B2 6 7 jjmit area=B2
IB1 0 5 pwl(0 0 5p IB1)
L1 a 1 2.082E-12
L2 1 4 2.06E-12
L3 4 6 2.067E-12
L4 6 q 2.075E-12
LP1 2 0 4.998E-13
LP2 7 0 5.011E-13
LB1 5 4 LB1
RB1 1 3 RB1
RB2 6 8 RB2
LRB1 3 0 LRB1
LRB2 8 0 LRB2
.ends
.ends
.ends