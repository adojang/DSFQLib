* JSIM deck file generated with TimEx
* === DEVICE-UNDER-TEST ===

* === SOURCE DEFINITION ===
.SUBCKT SOURCECELL  8 11
b1   1  2  jjmitll100 area=2.25
b2   3  4  jjmitll100 area=2.25
b3   5  6  jjmitll100 area=2.5
ib1  0  2  pwl(0 0 5p 275ua)
ib2  0  5  pwl(0 0 5p 175ua)
l1   8  7  1p
l2   7  0  3.9p
l3   7  1  0.6p
l4   2  3  1.1p
l5   3  5  4.5p
l6   5  11 2p
lp2  4  0  0.2p
lp3  6  0  0.2p
lrb1 9  2  1p
lrb2 10 4  1p
lrb3 12 6  1p
rb1  1  9  4.31
rb2  3  10 4.31
rb3  5  12 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS SOURCECELL
* === INPUT LOAD DEFINITION ===
.SUBCKT LOADINCELL  2 5
b1 1 6 jjmitll100 area=2.5
b2 4 8 jjmitll100 area=2.5
ib1 0 3 pwl(0 0 5p 350ua)
l1 2 1 2p
l2 1 3 2p
l3 3 4 2p
l4 4 5 2p
lb1 7 6 1p
lb2 9 8 1p
lp1 6 0 0.2p
lp2 8 0 0.2p
rb1 1 7 3.88
rb2 4 9 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS LOADINCELL
* === OUTPUT LOAD DEFINITION ===
.SUBCKT LOADOUTCELL  2 5
b1 1 6 jjmitll100 area=2.5
b2 4 8 jjmitll100 area=2.5
ib1 0 3 pwl(0 0 5p 350ua)
l1 2 1 2p
l2 1 3 2p
l3 3 4 2p
l4 4 5 2p
lb1 7 6 1p
lb2 9 8 1p
lp1 6 0 0.2p
lp2 8 0 0.2p
rb1 1 7 3.88
rb2 4 9 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS LOADOUTCELL
* === SINK DEFINITION ===
.SUBCKT SINKCELL  1
r1 1 0 2
.ENDS SINKCELL
* ===== MAIN =====
.param cval=600u
I_a 0 1000 pwl(0 0 
+500p 0 503p cval 505p 0 
+1000p 0 1003p cval 1005p 0)

*I_a 0 1000 pulse(0 600u 500p 2p 2p 1p 100p)
I_ext_clk 0 ext_clk pulse(0 600u 100p 2p 2p 1p 100p)

I_int_clk 0 int_clk pulse(0 600u 100p 2p 2p 1p 20p)
.tran 0.25p 1400p 0 0.01p

XSOURCEINa SOURCECELL 1000 2000
XLOADINa LOADINCELL 2000 A


XLOADOUTq LOADOUTCELL q 8000
XSINKOUTq SINKCELL 8000

XDFF1 LSmitll_DFF A ext_clk B
XNOT1 LSMITLL_NOT B int_clk D

*XSPLIT LSmitll_SPLIT int_clk clk1 clk2
*XJTL_Delay LSMITLL_JTL int_clk delay2
*XJTL_Delay2 LSMITLL_JTL delay2 delay3
*XJTL_Delay3 LSMITLL_JTL delay3 delay_clk

XNOT2 LSMITLL_NOT D int_clk F
XDFF2 LSmitll_DFF F ext_clk q

.subckt storage in out
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)



L1 in out 10p
RL out 1 0.5
BD 1 0 jjmit area=0.7
B1 out 0 jjmit area=1
RH out 0 4

.ends

.print v(B) v(D)
*.print i(L6.XSOURCEINa) i(I_ext_clk) i(L7.XDFF1) i(L12.XNOT1) i(L12.XNOT2) i(r1.XSINKOUTq) p(r1.XSINKOUTq)
*.print i(L6.XSOURCEINa) i(r1.XSINKOUTq)
*.print i(L4.XJTL_Delay3) i(L1.XNOT2) i(L12.XNOT2)


***************** NOT GATE *************************

*$Ports  a clk q
.subckt LSMITLL_NOT a clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=2.57
.param B3=1.07
.param B4=IC
.param B5=1.34
.param B6=3.03
.param B7=1.38
.param B8=0.8
.param B9=IC

.param IB1=BiasCoef*Ic0*B1
.param IB2=87u
.param IB3=257u
.param IB4=BiasCoef*Ic0*B4
.param IB5=BiasCoef*Ic0*B9

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9

.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet

.param RD=4
.param LRD=2p

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 7 8 jjmit area=B3
B4 13 14 jjmit area=B4
B5 17 18 jjmit area=B5
B6 10 11 jjmit area=B6
B7 20 18 jjmit area=B7
B8 18 19 jjmit area=B8
B9 21 22 jjmit area=B9

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 9 pwl(0 0 5p IB3)
IB4 0 15 pwl(0 0 5p IB4)
IB5 0 23 pwl(0 0 5p IB5)

LB1 3 1 LB1
LB2 6 4 LB2
LB3 8 9 LB3
LB4 13 15 LB4
LB5 21 23 LB5

L1 a 1 2.062E-12
L2 1 4 1.889E-12
L3 4 7 2.72E-12
L4 clk 13 2.057E-12
L5 13 16 1.029E-12
L6 16 17 1.241E-12
L7 16 12 1.973E-12
L8 10 12 1.003E-12
L9 10 8 7.524E-12
L10 8 20 1.234E-12
L11 18 21 2.607E-12
L12 21 q 2.062E-12

LP1 2 0 5.271E-13
LP2 5 0 5.237E-13
LP4 14 0 4.759E-13
LP6 11 0 5.021E-13
LP8 19 0 6.33E-13
LP9 22 0 4.749E-13

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 5 LRB2
RB3 7 107 RB3
LRB3 107 8 LRB3
RB4 13 113 RB4
LRB4 113 0 LRB4
RB5 17 117 RB5
LRB5 117 18 LRB5
RB6 10 110 RB6
LRB6 110 0 LRB6
RB7 20 120 RB7
LRB7 120 18 LRB7
RB8 18 118 RB8
LRB8 118 0 LRB8
RB9 21 121 RB9
LRB9 121 0 LRB9
LRD 12 112 LRD
RD 112 0 RD
.ends

***************** DFF CELL *************************


*$Ports		a		clk		q
.subckt LSmitll_DFF	  a	clk q	
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.70

.param B1=2.5
.param B2=1.61
.param B3=1.54
.param B4=1.69
.param B5=1.38
.param B6=2.5
.param B7=2.5

.param IB1=175u     
.param IB2=173u      
.param IB3=175u            
.param IB4=175u        

.param L1=Phi0/(4*IC*Ic0)               
.param L2=Phi0/(2*B1*Ic0)         
.param L3=Phi0/(B3*Ic0)       
.param L4=Phi0/(2*B6*Ic0)      
.param L5=Phi0/(4*IC*Ic0)     
.param L6=Phi0/(2*B4*Ic0)       
.param L7=Phi0/(4*B7*Ic0)         
.param LB1=LB            
.param LB2=LB           
.param LB3=LB           
.param LB4=LB        
.param LP1=LP         
.param LP3=LP          
.param LP4=LP         
.param LP6=LP          
.param LP7=LP          
.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2       
.param RB3=B0Rs/B3          
.param RB4=B0Rs/B4         
.param RB5=B0Rs/B5         
.param RB6=B0Rs/B6          
.param RB7=B0Rs/B7
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 5 6 jjmit area=B3
B4 8 9 jjmit area=B4
B5 10 8 jjmit area=B5
B6 11 12 jjmit area=B6
B7 14 15 jjmit area=B7

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 13 pwl(0 0 5p IB3)
IB4 0 16 pwl(0 0 5p IB4)

LB1 3 1 LB1
LB2 7 5 LB2
LB3 11 13 LB3
LB4 16 14 LB4

L1 a 1 2.059E-12
L2 1 4 4.123E-12
L3 5 8 6.873E-12
L4 10 11 5.195E-12
L5 clk 11 2.071E-12
L6 8 14 3.287E-12
L7 14 q 2.066E-12

LP1 2 0 5.042E-13    
LP3 6 0 5.799E-13    
LP4 9 0 5.733E-13    
LP6 12 0 4.605E-13    
LP7 15 0 4.961E-13    

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 5 LRB2
RB3 5 105 RB3
LRB3 105 0 LRB3
RB4 8 108 RB4
LRB4 108 0 LRB4
RB5 10 110 RB5
LRB5 110 8 LRB5
RB6 11 111 RB6
LRB6 111 0 LRB6
RB7 14 114 RB7
LRB7 114 0 LRB7
.ends



********************** JTL *****************************
*$Ports 			a q
.subckt LSMITLL_JTL a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=IC
.param IB1=(B1+B2)*Ic0*BiasCoef
.param LB1=LB
.param L1=Phi0/(4*B1*Ic0)
.param L2=Phi0/(4*B1*Ic0)
.param L3=Phi0/(4*B1*Ic0)
.param L4=Phi0/(4*B2*Ic0)
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP

B1 1 2 jjmit area=B1
B2 6 7 jjmit area=B2
IB1 0 5 pwl(0 0 5p IB1)
L1 a 1 2.082E-12
L2 1 4 2.06E-12
L3 4 6 2.067E-12
L4 6 q 2.075E-12
LP1 2 0 4.998E-13
LP2 7 0 5.011E-13
LB1 5 4 LB1
RB1 1 3 RB1
RB2 6 8 RB2
LRB1 3 0 LRB1
LRB2 8 0 LRB2
.ENDS

.end
