* A Generic flipflopflop for simulating Logic Gates
* Copyright (c) 2022-2024 Adriaan van Wijk, Stellenbosch University
*


.tran 0.25p 1000p 0 0.25p



*VsrcA 1 0 pwl(0 0 50p 0 51p 600u 52p 0)

.model J0 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)

.model J1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=132uA)

.model J70 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=70uA)

.model J141 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=141uA)

.model J350 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=350uA)

.model J2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=513uA)

I0 0 1 pwl(0 0 5p 100u)



I1 0 3 pwl(0 0 5p 100u)
I2 0 4 pwl(0 0 5p 411u)
I3 0 7 pwl(0 0 5p 100u)
Ib61 0 100 pwl(0 0 5p 263u)
Ib62 0 flop_S pwl(0 0 5p 263u)


L0 1 2 8p
L1 3 4 4p
L2 4 5 0.973p
L3 flop_S 6 3p
L4 7 8 25p
L5 8 F 4p
L6 9 101 4p
L7 5 100 4p
L8 5 flop_S 4p


B0 2 3 J0
Rb0 2 33 1
Lb0 33 3 0.7p

B1 3 0 J1
Rb1 3 30 1
Lb1 30 0 0.7p

B2 4 0 0 J2
Rb2 4 99 1
Lb2 99 0 0.7p

B3 6 7 J0
Rb3 6 77 1
Lb3 77 7 0.7p

B4 7 0 J141
Rb4 7 70 1
Lb4 70 0 0.7p

B5 8 0 J141
Rb5 8 88 1
Lb5 88 0 0.7p

B6 8 9 J0
Rb6 8 900 1
Lb6 900 9 1p

B61 100 0 J350
R61b 100 611 1
L61b 611 0 1p

B62 flop_S 0 J350
R62b flop_S 612 1
L62b 612 0 1p




Rs F 0 2

*Testing Dynamic Hold times

Lp 100 101 10p
Rl 101 102 0.5
Bd 102 0 J70
Bj 101 0 J0
Rh 101 0 4


.print v(1) v(3) v(5) v(flop_S) v(101) v(8) v(Rs)
*.print p(B0) p(B1) p(B2) p(B3) p(B5)

.end


josim -o ./test.csv ./test.cir -V 1
josim-plot.py ./test.csv -t stacked
