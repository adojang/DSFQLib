* JSIM deck file generated with TimEx
* This testbench uses the AW_AND_base.cir file

* === SOURCE DEFINITION ===
.SUBCKT SOURCECELL  8 11
b1   1  2  jjmitll100 area=2.25
b2   3  4  jjmitll100 area=2.25
b3   5  6  jjmitll100 area=2.5
ib1  0  2  pwl(0 0 5p 275ua)
ib2  0  5  pwl(0 0 5p 175ua)
l1   8  7  1p
l2   7  0  3.9p
l3   7  1  0.6p
l4   2  3  1.1p
l5   3  5  4.5p
l6   5  11 2p
lp2  4  0  0.2p
lp3  6  0  0.2p
lrb1 9  2  1p
lrb2 10 4  1p
lrb3 12 6  1p
rb1  1  9  4.31
rb2  3  10 4.31
rb3  5  12 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS SOURCECELL
* === INPUT LOAD DEFINITION ===
.SUBCKT LOADINCELL  2 5
b1 1 6 jjmitll100 area=2.5
b2 4 8 jjmitll100 area=2.5
ib1 0 3 pwl(0 0 5p 350ua)
l1 2 1 2p
l2 1 3 2p
l3 3 4 2p
l4 4 5 2p
lb1 7 6 1p
lb2 9 8 1p
lp1 6 0 0.2p
lp2 8 0 0.2p
rb1 1 7 3.88
rb2 4 9 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS LOADINCELL
* === OUTPUT LOAD DEFINITION ===
.SUBCKT LOADOUTCELL  2 5
b1 1 6 jjmitll100 area=2.5
b2 4 8 jjmitll100 area=2.5
ib1 0 3 pwl(0 0 5p 350ua)
l1 2 1 2p
l2 1 3 2p
l3 3 4 2p
l4 4 5 2p
lb1 7 6 1p
lb2 9 8 1p
lp1 6 0 0.2p
lp2 8 0 0.2p
rb1 1 7 3.88
rb2 4 9 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS LOADOUTCELL
* === SINK DEFINITION ===
.SUBCKT SINKCELL  1
r1 1 0 2
.ENDS SINKCELL
* ===== MAIN =====
.param cval=600u

I_a 0 1000 pwl(0 0 
+100p 0 103p cval 105p 0
+300p 0 303p cval 305p 0
+350p 0 353p cval 355p 0
+400p 0 403p cval 405p 0
+450p 0 453p cval 455p 0
+500p 0 503p cval 505p 0
+710p 0 713p cval 715p 0
+820p 0 823p cval 825p 0
+850p 0 853p cval 855p 0)

I_b 0 4000 pwl(0 0 
+200p 0 203p cval 205p 0
+300p 0 303p cval 305p 0
+350p 0 353p cval 355p 0
+405p 0 408p cval 410p 0
+460p 0 463p cval 465p 0
+515p 0 518p cval 520p 0
+710p 0 713p cval 715p 0
+820p 0 823p cval 825p 0
+850p 0 853p cval 855p 0)


XSOURCEINa SOURCECELL 1000 2000
XLOADINa LOADINCELL 2000 A

XSOURCEINb SOURCECELL 4000 5000
XLOADINb LOADINCELL 5000 B
XLOADOUTq LOADOUTCELL q 8000
XSINKOUTq SINKCELL 8000

*XDUT DSFQ_AND A B q

.tran 0.25p 600p 0 0.01p
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)



*$Ports    A B q
*.subckt DSFQ_AND A B q

* The throughput for this logic cell is approximately 5ps with zero skew applied.
* The skew tolerance can be adjusted using the following formula:
* RHold = a * (16.666 * t_hold)^b
* Where a = 3.572e-10
* and   b = -1.023


* 				*(*************************** VERSION 1.3 of the AND GATE STARTS HERE *****************************************)

.param  b1  	=	 	 3.23682804e-01
.param  b2  	=	 	 5.95629005e-01
.param 	b3 		= 		 b1
.param 	b4 		= 		 b2
.param  b5  	=	 	 6.21776921e-01
.param  i1  	=	 	 3.00270413e-05
.param  l1  	=	 	 5.22896652e-12
.param 	l2 		= 		 l1
.param  l3  	=	 	 1.73951938e-12
.param  lp1  	=	 	 9.19415844e-14
.param  lrb1  	=	 	 4.30836486e-12
.param  lrb2  	=	 	 7.59006914e-12
.param  lrb3  	=	 	 5.78336737e-12
.param  lrb4  	=	 	 1.55573615e-12
.param  lrb5  	=	 	 1.06776433e-12
.param  ra  	=	 	 2.41454521e+00
.param  rb1  	=	 	 3.27679568e+00
.param  rb2  	=	 	 4.66908026e+00
.param 	rb3 	= 		 rb1
.param 	rb4 	= 		 rb2
.param  rb5  	=	 	 7.26286283e+00

* Back Annotated .cir file from KiCad
b1   	4   	5   	 jjmit area=b1
b2   	6   	7   	 jjmit area=b2
b3   	4   	8   	 jjmit area=b3
b4   	6   	4   	 jjmit area=b4
b5   	4   	9   	 jjmit area=b5
i1   	0   	4   	pwl(0   	0   	5p   	i1)
l1   	a   	5   	 l1
l2   	b   	7   	 l1
l3   	4   	q   	 l3
lp1   	9   	0   	 lp1
lrb1   	10   	4   	 lrb1
lrb2   	11   	6   	 lrb2
lrb3   	12   	4   	 lrb1
lrb4   	13   	6   	 lrb2
lrb5   	14   	0   	 lrb5
r1   	8   	5   	 rA
r2   	4   	7   	 rA
r3   	5   	4   	 rA
r4   	7   	6   	 rA
rb1   	5   	10   	 rb1
rb2   	7   	11   	 rb2
rb3   	8   	12   	 rb3
rb4   	4   	13   	 rb4
rb5   	4   	14   	 rb5


*.print v(L4.XLOADINa) v(r1.XSINKOUTq) v(L4.XLOADINb) p(B5.XDUT)
.print p(B5)

.end