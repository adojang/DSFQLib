.subckt master A B C Q
.param R1   =   5

* xtest1 one A B Q1
Lxtest1_1 A A_one 0
Lxtest2_2 B B_one 0
Lxtest3_3 Q Q1_one 0

* xtest2 two Q1 C Q
Lxtest1_1 Q1 A_two 0
Lxtest2_2 C B_two 0
Lxtest3_3 Q Q_two 0

* .subckt one A B Q
.param Lp   =   5
.param b1   =   1
.param i1   =   1
L1 A_one AA_one Lp
L2 B_one BB_one 15
R1 A_one 0 20
b1   	30_one   	10_one   	 jjmit area=b1_one
i1   	0   	30_one   	pwl(0   	0   	5p   	i1_one)
* xtest3 three AA BB
Lxtest3_1 AA_one Ax_three_one 0
Lxtest3_2 BB_one Bx_three_one 0
* .subckt three Ax Bx
.param Lp_three_one   =   5
.param b1_three_one   =   1
.param i1_three_one   =   1
L1 25_three_one Ax_three_one Lp_three_one
L2 15_three_one Bx_three_one 15
R1 Bx_three_one 0 20
b1   	30_three_one   	10_three_one   	 jjmit area=b1_three_one
i1   	0   	30_three_one   	pwl(0   	0   	5p   	i1_three_one)
* .ends
* .ends


*.subckt two A B Q
.param Lp_two   =   5
.param b1_two   =   1
.param i1_two   =   1
L1 0 A_two Lp_two
L2 15_two B_two 15
R1 15_two Q_two 20
b1   	30_two   	10_two   	 jjmit area=b1_two
i1   	0   	30_two   	pwl(0   	0   	5p   	i1_two)
*.ends
.ends