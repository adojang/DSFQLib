*.include LSmitll_JTL_v2p1_optimized.cir
*Comment the line above to see results. Ideally it should be included, but because it is included \
*In the main .cir file, this causes an error. This is a temporary solution meanwhile...

.include AW_mitll_OR_optimized.cir
.include AW_mitll_AND_optimized.cir
*.include LSmitll_SPLIT_v2p1_optimized.cir
.include LSmitll_NOT_v2p1_optimized.cir

*Propagation Delay Times:
*XSPLIT -   12ps
*XMRG   -   9ps
*XOR    -   16ps
*Total =    48ps (longest path xyz)

.subckt DSFQ_2_1_MUX A0 B0 S0 QQ
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)

XSPLITA LSMITLL_SPLIT A0 A1 CLK
XSPLITS LSMITLL_SPLIT S0 S1 B2

XDELAYB  LSMITLL_JTL B0 B1

XNOT    LSMITLL_NOT   S1 CLK A2
XAND1   DSFQ_AND   A1 A2 Q1
XAND2   DSFQ_AND   B1 B2 Q2
XOR     DSFQ_OR    Q1 Q2 QQ
.ends