.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_SFQDC_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include AW_mitll_DSFQ_NOT.cir

.tran 0.025p 400p 0
.param cval= 600u

I_A0 0 xa pwl(0 0 100p 0 103p cval 105p 0 200p 0 203p 0 205p    0 300p 0 303p cval 305p 0) 
I_B0 0 xb pwl(0 0 150p 0 153p cval 155p 0 107p 0 110p 0 112p 0 200p 0 203p cval 205p 0 300p 0 303p    0 305p 0)
I_C0 0 xc pwl(0 0 100p 0 103p 0 105p 0 108p 0 111p 0 113p 0 200p 0 203p 0 205p 0 300p 0 303p    0 305p 0)

*Expected Outputs: 0 1 0

XDCSFQA LSmitll_DCSFQ xa xa1 
XDCSFQB LSmitll_DCSFQ xb xb1
XDCSFQC LSmitll_DCSFQ xc xc1 

XJTLA LSMITLL_JTL xa1 A
XJTLB LSMITLL_JTL xb1 B
XJTLC LSMITLL_JTL xc1 C

XNOT MASTER A B C Q

XLOAD LSMITLL_JTL q qq

Rsink qq 0 2

.print  p(A) p(CLK1.XNOT) p(Q)



******* INCLUDED FILES *******


*.subckt master a b c q
.param lad  	=	 	    5

xtest1 one a b q1
xtest2 two q1 c q

*.subckt one am bm q1m
l_connect_0 xaa xaa 0

l_connect_1 xbb xbb 0

l1 am xaa 5
r1 xbb bm 5
c1 xbb qm1
xtest3 three saa_three_one sbb_three_one


*.subckt three saa sbb
l_connect_0_three xrr_three xrr_three 0

l_connect_1_three xyy_three xyy_three 0

l1_three saa_three fr1_three 55
lr_three fr1_three xrr_three 553
lk_three xyy_three sbb_three 33

xrinox rhino oupa_rhino_three_one hannes_rhino_three_one

*.subckt rhino oupa hannes
.param opsies_rhino_three = 55
.param katjie_rhino_three = 767
r1_rhino_three oupa_rhino_three hannes_rhino_three opsies_rhino_three
r2_rhino_three hannes_rhino_three 0 katjie_rhino_three
*.ends


*.ends


*.ends

*.ends

*.ends


*.subckt two q1m cm q
l1_two q1m_two cm_two 5
r1_two q1_two 0 5
c1_two q11_two q_two *.ends_two




*.ends