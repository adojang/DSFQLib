.title KiCad schematic
R2 /22 /20 Resistor
B8 /40 /31 jjmit
L6 /40 Q Inductor
LP5 /31 GND Inductor
LP4 /24 GND Inductor
B9 /24 /22 jjmit
LC1 /10a /10b Inductor
B3 /3 /10a jjmit
B4 /5 /3 jjmit
LP1 /5 GND Inductor
B2 /4 /2 jjmit
B1 /3 /1 jjmit
L1 A /1 Inductor
L2 B /2 Inductor
LC2 /10b /10c Inductor
LBIAS1 /biasa /10b Inductor
RBIAS1 /biasa bias Resistor
L3 /10b /30 Inductor
LP2 /6 GND Inductor
LC3 /30 /40 Inductor
L4 /30 /20 Inductor
R1 /21 /20 Resistor
B7 /24a /20 jjmit
LR1 /21 /24 Inductor
LB7 /24a /24 Inductor
B5 /4 /10c jjmit
B6 /6 /4 jjmit
LP3 /24 GND Inductor
.end
