* DSFQ Self clocked Multiplexor
* Author: Adriaan van Wijk
* Version: 1.0
* Last modification date: 21 June 2022
* Last modification by: Adriaan van Wijk
* This testbench uses cells from LS's library of RSFQ cells. This was the version that was tested for layout.

.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
*JTL Conflicts with what is already in the MUX cell. It is a Bug(?).
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include cells\AW_2_1_MUX.cir

*SPLIT Conflicts with what is already in the MUX Cell. It is a Bug.
.include cells\LSmitll_SPLIT_v2p1_optimized.cir 

.param cval=600u

********************************************* THROUGHPUT TIMES ROUGHLY ********************************************
*i0 output time: 112ps two levels. Inputs A-A
*i1 output time: 90ps - two levels. Inputs B-A
*i2 output time: 90ps - Inputs A-B
*i3 output time: 70ps - Inputs B-B

*Everything is able to output. The problem lies in the stacking of timing errors between the A and B inputs since the internals are not balanced.
*Suggest a MUX redesign to balance things properly, and a better overview.
********************************************* THROUGHPUT TIMES ROUGHLY ********************************************

* I_i0 0 i_i0 pwl(0 0 100p 0 103p 0 105p 0 200p 0 203p 0 205p 0 300p 0 303p 0 305p 0 400p 0 403p 0 405p 0 500p 0 503p cval 505p 0)
* I_i1 0 i_i1 pwl(0 0 100p 0 103p 0 105p 0 200p 0 203p 0 205p 0 300p 0 303p 0 305p 0 400p 0 403p 0 405p 0 500p 0 503p 0 505p 0)
* I_i2 0 i_i2 pwl(0 0 100p 0 103p 0 105p 0 200p 0 203p 0 205p 0 300p 0 303p 0 305p 0 400p 0 403p 0 405p 0 500p 0 503p 0 505p 0)
* I_i3 0 i_i3 pwl(0 0 100p 0 103p cval 105p 0 200p 0 203p 0 205p 0 300p 0 303p 0 305p 0 400p 0 403p 0 405p 0 500p 0 503p 0 505p 0)

* I_s0 0 i_s0 pwl(0 0 130p 0 133p cval 135p 0 200p 0 203p 0 205p 0 320p 0 323p 0 325p 0 420p 0 423p 0 425p 0 500p 0 503p 0 505p 0)
* I_s1 0 i_s1 pwl(0 0 100p 0 103p cval 105p 0 200p 0 203p 0 205p 0 300p 0 303p 0 305p 0 400p 0 403p 0 405p 0 500p 0 503p 0 505p 0)


I_i0 0 i_i0 pwl(0 0 100p 0 103p cval 105p 0 200p 0 203p 0 205p 0 300p 0 303p 0 305p 0 400p 0 403p 0 405p 0 500p 0 503p 0 505p 0)
I_i1 0 i_i1 pwl(0 0 100p 0 103p 0 105p 0 200p 0 203p cval 205p 0 300p 0 303p 0 305p 0 400p 0 403p 0 405p 0 500p 0 503p 0 505p 0)
I_i2 0 i_i2 pwl(0 0 100p 0 103p 0 105p 0 200p 0 203p 0 205p 0 300p 0 303p cval 305p 0 400p 0 403p 0 405p 0 500p 0 503p 0 505p 0)
I_i3 0 i_i3 pwl(0 0 100p 0 103p 0 105p 0 200p 0 203p 0 205p 0 300p 0 303p 0 305p 0 400p 0 403p cval 405p 0 500p 0 503p 0 505p 0)

I_s0 0 i_s0 pwl(0 0 100p 0 103p 0 105p 0 200p 0 203p 0 205p 0 320p 0 323p cval 325p 0 420p 0 423p cval 425p 0 500p 0 503p 0 505p 0)
I_s1 0 i_s1 pwl(0 0 100p 0 103p 0 105p 0 200p 0 203p cval 205p 0 300p 0 303p 0 305p 0 400p 0 403p cval 405p 0 500p 0 503p 0 505p 0)

*S0 must be delayed by ~30ps for things to work properly. This realtes to Q2's MUX.


* I_i2 0 i_i2 pwl(0 0 300p 0 303p cval 305p 0)
* I_s0 0 i_s0 pwl(0 0 300p 0 303p cval 305p 0)
* I_s1 0 i_s1 pwl(0 0 300p 0 303p 0 305p 0)

*Design a test which outputs i0 i1 i2 i3 sucessfully.


.tran 0.25p 600p 0 0.01p
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)

Xsrc_i0 LSmitll_DCSFQ i_i0 src_i0
Xsrc_i1 LSmitll_DCSFQ i_i1 src_i1
Xsrc_i2 LSmitll_DCSFQ i_i2 src_i2
Xsrc_i3 LSmitll_DCSFQ i_i3 src_i3
Xsrc_s0 LSmitll_DCSFQ i_s0 src_s0
Xsrc_s1 LSmitll_DCSFQ i_s1 src_s1


Xload_i0 LSMITLL_JTL src_i0 i0
Xload_i1 LSMITLL_JTL src_i1 i1
Xload_i2 LSMITLL_JTL src_i2 i2
Xload_i3 LSMITLL_JTL src_i3 i3
Xload_s0 LSMITLL_JTL src_s0 S0
Xload_s1 LSMITLL_JTL src_s1 S1

XSPLITS LSMITLL_SPLIT S1 S1A S1B


XMUXA   DSFQ_2_1_MUX i0 i1 S1A Q1
XMUXB   DSFQ_2_1_MUX i2 i3 S1B Q2
XMUXC   DSFQ_2_1_MUX Q1 Q2 S0 QQ

Xloadout_s0 LSMITLL_JTL QQ Qload
R_out Qload 0 2




*I might need to insert a small JTL type element on A1 and B1 inside the 2:1 MUX for stability. Might need to do the same for Q1 and Q2 in teh 2-1 MUX.

*.print v(i2) v(Q2)  p(A1.XMUXB) v(A_clk.XMUXB) v(S1.XMUXB) v(A2.XMUXB) p(A2.XMUXB) p(Q1.XMUXB)



*1 2 3 4 Test Pattern Print Confirmation
.print v(i0) v(i2) v(i1) v(i3) v(Q1) v(Q2) v(s1) v(s0)  v(QQ)


*Test Confirmation:

* 100 ps
* i0 high i2 high i3 high
* s1 high s1 high

* Q1 should be i1 =low
* Q2 should be i3 = high
* QQ should be Q1 = low
* True? YES.

* 200 ps
* i0 low i1 high i2 low i3 low
* s1 high s0 low
* Q1 should be i1 = high
* Q2 should be i3 = low
* QQ should be Q1 = high
* True? FALSE. Q1 does not switch. Why?



*Time 3 troubleshooting
*.print v(i2) v(s1) p(Q1) p(Q2) p(QQ)  p(S1.XMUXB) p(CLK_BOOST.XMUXB) p(A2.XMUXB)

* ON: i0 i2 i3
* Selected: (0 - A, 1 - B) S1 = 1 therefore B therefore i1 and i3.
* i3 is ON therefore Q2 is ON i1 is off therefore Q1 is OFF
* Q1 OFF Q2 ON Select line is 0 therefore output OFF
*Output QQ should be LOW
* PASS


* At time 200ps
* i1 = ON all else is off
* S1 is on, therefore B input high
* i1 = 1 therefore Q1 =1
* i3 = = therefore Q2 =0
* S0 = 0 therefore A input therefore Q1.
*Output QQ should be HIGH
* PASS

* at time 300ps
* i2 = HIGH all else LOW
* S1 = LOW therefore A input therefore i2 input
* We expect Q1 - LOW and Q2 HIGH
* Q2 should be HIGH but is not HIGH. Inverting clk bug.
* S0 HIGH so B input select Q2
* OUTPUT SHOULD BE HIGH FOR QQ BUT IS NOTT.

* ===============================
* The problem lies in the OR Gate I think. Something is causing the NOT gate to have low outputs. I think its the inputs.
* PRoblem defs lies in teh OR gate. We have a: HIGH, Semi-low combo that outputs a HALF high. Very broken indeed.

*.print v(i0) v(S1.XMUXA) v(CLK.XMUXA) v(A2.XMUXA) v(Q1.XMUXA) v(Q2.XMUXA) v(Q1)
*.print v(S0) v(S1) v(AA)


.end