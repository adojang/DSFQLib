* DSFQ Self clocked Multiplexor
* Author: Adriaan van Wijk
* Version: 1.0
* Last modification date: 21 June 2022
* Last modification by: Adriaan van Wijk
* This testbench uses cells from LS's library of RSFQ cells. This was the version that was tested for layout.

.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include cells\LSmitll_SPLIT_v2p1_optimized.cir
.include AW_mitll_DSFQ_AND.cir
.include AW_mitll_DSFQ_OR.cir
.include AW_mitll_DSFQ_XOR.cir
.include cells\LSmitll_BUFF_v2p1_optimized.cir
.param cval=600u

I_a0 0 I_a0 pwl(0 0 100p 0 103p 0 105p 0        200p 0 203p 0 205p 0         300p 0 303p 0 305p 0        400p 0 403p cval 405p 0        500p 0 503p cval 505p 0         600p 0 603p cval 605p 0         700p 0 703p cval 705p 0)
I_b0 0 I_b0 pwl(0 0 100p 0 103p 0 105p 0     200p 0 203p cval 205p 0      300p 0 303p cval 305p 0     400p 0 403p 0 405p 0           500p 0 503p 0 505p 0            600p 0 603p cval 605p 0         700p 0 703p cval 705p 0)
I_ci 0 I_ci pwl(0 0 100p 0 103p cval 105p 0     200p 0 203p 0 205p 0         300p 0 303p cval 305p 0     400p 0 403p 0 405p 0           500p 0 503p cval 505p 0         600p 0 603p 0 605p 0            700p 0 703p cval 705p 0)
I_s0 0 I_s0 pwl(0 0 170p 0 173p cval 175p 0     270p 0 273p cval 275p 0      370p 0 373p 0 375p 0        470p 0 473p cval 475p 0        570p 0 573p 0 575p 0            670p 0 673p 0 675p 0            770p 0 773p cval 775p 0)
I_z0 0 I_z0 pwl(0 0 100p 0 103p 0 105p 0        200p 0 203p 0 205p 0         300p 0 303p cval 305p 0     400p 0 403p 0 405p 0           500p 0 503p cval 505p 0         600p 0 603p cval 605p 0         700p 0 703p cval 705p 0)
*S = 0 - Select A
*S = 1 - Select B

* A   0 0 0 1 1 1 1
* B   0 1 1 0 0 1 1
* Ci  1 0 1 0 1 0 1
* S   1 1 0 1 0 0 1
* Cot 0 0 1 0 1 1 1


.tran 0.25p 800p 0 0.05p

Xsrc_a0 LSmitll_DCSFQ i_a0 src_a0
Xsrc_b0 LSmitll_DCSFQ i_b0 src_b0
Xsrc_ci LSmitll_DCSFQ i_ci src_ci
Xsrc_s0 LSmitll_DCSFQ i_s0 src_s0
Xsrc_z0 LSmitll_DCSFQ i_z0 src_z0

Xload_a0 LSMITLL_JTL src_a0 A0
Xload_b0 LSMITLL_JTL src_b0 B0
Xload_c0 LSMITLL_JTL src_ci Cin
Xload_s0 LSMITLL_JTL src_s0 S_BASE
Xload_z0 LSMITLL_JTL src_z0 Carry_BASE

*For Reference to confirm it is working correctly.
R_QS S_BASE 0 4
R_Cout Carry_BASE 0 4

XSPTA LSMITLL_SPLIT A0 A11 A22
XSPTB LSMITLL_SPLIT B0 B11 B22
XJTLA1 LSMITLL_JTL  A11 A1
XJTLB1 LSMITLL_JTL  B11 B1
XJTLA2 LSMITLL_JTL  A22 A2
XJTLB2 LSMITLL_JTL  B22 B2

XXOR3 DSFQ_XOR Cin 0 C0
XSPTC LSMITLL_SPLIT C0 C11 C22

XJTLC1 LSMITLL_JTL  C11 C101
XJTLC101 LSMITLL_JTL  C101 C102
XJTLC102 LSMITLL_JTL  C102 C103
XJTLC103 LSMITLL_JTL  C103 C1

XJTLC2 LSMITLL_JTL  C22 C201
XJTLC201 LSMITLL_JTL  C201 C202
XJTLC202 LSMITLL_JTL  C202 C203
XJTLC203 LSMITLL_JTL  C203 C2

XXOR1 DSFQ_XOR A1 B1 XOR0
XJTLXOR LSMITLL_JTL  XOR0 XOR1
XSPTD LSMITLL_SPLIT XOR1 XOR1aa XOR1bb
XJTLXOR1a LSMITLL_JTL  XOR1aa XOR1a
XJTLXOR1b LSMITLL_JTL  XOR1bb XOR1b

XXOR2 DSFQ_XOR C1 XOR1a S

XAND1 DSFQ_AND A2 B2 AND11
XAND2 DSFQ_AND XOR1b C2 AND22
XJTLAND1 LSMITLL_JTL  AND11 AND1
XJTLAND2 LSMITLL_JTL  AND22 AND2

XOR DSFQ_OR AND1 AND2 Cout
.print p(S_BASE) p(Carry_BASE) p(Sout)  p(CarryOut)
*  .print p(S_BASE) p(Carry_BASE) p(S)  p(Cout) p(AND1) p(XOR1b) p(AND2) p(C2) p(XOR1b) p(C1)

XCOUT LSMITLL_JTL Cout Carryout
R_Carry Carryout 0 2
XLOAD LSMITLL_JTL S Sout
R_out Sout 0 2

.end