.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_SFQDC_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include AW_mitll_DSFQ_AND.cir

.tran 0.015p 500p 0
.param cval= 600u

*15ps skew with 2e-12 input.
I_A0 0 xa pwl(0 0 100p 0 103p cval 105p 0 200p 0 203p 0 205p 0 300p 0 303p cval 305p 0   400p 0 403p cval 405p 0) 
I_B0 0 xb pwl(0 0 100p 0 103p 0 105p 0 200p 0 203p cval 205p 0 300p 0 303p cval 305p 0      410p 0 413p cval 415p 0)
* I_A1 0 xc pwl(0 0 100p 0 103p cval 105p 0 200p 0 203p 0 205p 0) 
* I_B1 0 xd pwl(0 0 100p 0 103p cval 105p 0 213p cval 216p 0 218p 0)

*A   1 1
*B   0 1
*Q   0 1

XDCSFQA LSmitll_DCSFQ xa xa1 
XDCSFQB LSmitll_DCSFQ xb xb1

XJTLA LSMITLL_JTL xa1 A
XJTLB LSMITLL_JTL xb1 B

XDUT DSFQ_AND A B q

XLOAD LSMITLL_JTL q qq
Rsink qq 0 2

.print p(A) p(B) p(Q)