* A Generic DSFQ AND Gate for use in simulating Logic Gates
* Copyright (q) 2022-2024 Adriaan van Wijk, Stellenbosch University
* Based on the design by Rylov [2019]
*
* This gate is not meant to be directly attached to PTLs as it does not support integrated PTL ports.
* Version 1.0

*$Ports 		 A B q
.subckt DSFQ_AND A B q

.param main=0.84
.param secondary=0.60
.param third=1.68
.param pInduc = 1p
.param retentionResistor=4

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)

L1 A 1 12p
L2 B 4 12p
RD1 1 2 0.67
RD2 4 5 0.67

BD1 2 q jjmit area=secondary
RDp1 2 14 2.8
Ld1 14 q pInduc

BD2 5 q jjmit area=secondary
RDp2 5 15 2.8
Ld2 15 q pInduc

Rh1 1 q retentionResistor

B1 1 q jjmit area=main
Rb1 1 10 2.37
Lb1 10 q pInduc

Rh2 4 q retentionResistor

B2 4 q jjmit area=main
Rb2 4 11 2.37
Lb2 11 q pInduc

B3 0 q jjmit area=third
Rb3 q 13 1.67
Lb3 13 0 pInduc

Ibias 0 q dc 70u
.ends