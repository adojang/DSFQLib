.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_SFQDC_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include translated_shunt.cir
.tran 0.025p 250p 0
.param cval= 600u
I_A0 0 xa pwl(0 0 100p 0 103p cval 105p 0 200p 0 203p 0 205p 0) 
I_B0 0 xb pwl(0 0 122p 0 125p 0 127p 0 200p 0 203p 0 205p 0)
XDCSFQA LSmitll_DCSFQ xa xa1 
XDCSFQB LSmitll_DCSFQ xb xb1
XJTLA LSMITLL_JTL xa1 A
XJTLB LSMITLL_JTL xb1 B
XDUT RYLOV A B q
XLOAD LSMITLL_JTL q qq
Rsink qq 0 2
.print i(L1.XDUT)
.subckt RYLOV a b q
.param 	b1  	= 0.84
.param 	b2  	= 0.84
.param 	b3  	= 0.60
.param 	b4  	= 0.60
.param 	b5  	= 1.68
.param 	i1  	= 70u
.param l1 = 12.0p
.param l2 = 12.0p
.param 	l3  	= 2p
.param lp1      = 0.2p
.param 	lrb5  	= 2.3071p
.param 	r1  	= 4
.param 	r2  	= 4
.param 	r3  	= 0.68
.param 	r4  	= 0.68
.param 	rb5  	= 4.0833

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
* Back Annotated .cir file from KiCad
b1   	10   	39   	 jjmit area=b1
b2   	30   	20   	 jjmit area=b2
b3   	12   	39   	 jjmit area=b3
b4   	30   	22   	 jjmit area=b4
b5   	31   	30   	 jjmit area=b5
i1   	0   	30   	pwl(0   	0   	5p   	i1)
l1   	a   	10   	 l1
l2   	b   	20   	 l2
l3   	30   	q   	 l3
lp1   	31   	0   	 lp1
lrb5   	32   	0   	 lrb5
r1   	10   	39   	 r1

lmeasure      39      30      0

r2   	20   	30   	 r2
r3   	12   	10   	 r3
r4   	22   	20   	 r4
rb5   	30   	32   	 rb5
.ends
