* DC Pulse Generator
* Copyright (c) 2022-2024 Adriaan van Wijk, Stellenbosch University
*
* This pulse generator uses a DC current source to generate a SFQ pulse. The LSmitll DC to SFQ cell is used.

.tran 0.25p 200p 0 0.025p

.model J0 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=650uA)

.model J1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=132uA)

.model J2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=513uA)

I0 0 1 pwl(0 0 5p 650u)
I1 0 6 pwl(0 0 5p 100u)
I2 0 7 pwl(0 0 5p 411u)

L1 6 7 4p
L2 7 8 0.973p

XSFQ LSmitll_DCSFQ 4 6

B0 	2 4 J0
Rb0 2 2x 1
Lb0 2x 4 1p

B1 6 0 J1
Rb1 6 6x 1
Lb1 6x 0 0.7p

B2 7 0 0 J2
Rb2 7 7x 1
Lb2 7x 0 0.7p

*These values were tuned, not calculated.
LI 1 2 300p
RI 1 0 16



.print v(1) v(6) v(7)
*.print p(1) p(6) p(7)

*===== DC to SFQ Source =======
*$Ports 			a q
.subckt LSmitll_DCSFQ a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

.param B0=1.0
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LB=2p
.param LP=0.2p

.param B1=2.25
.param B2=2.25
.param B3=2.5
.param L1=1p
.param L2=3.9p
.param L3=0.6p
.param L4=1.1p
.param L5=4.5p
.param L6=2p
.param IB1=275u
.param IB2=175u
.param LB1=LB
.param LB2=LB
.param LP2=LP
.param LP3=LP
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet

B1 2 3 jjmit area=B1
B2 5 6 jjmit area=B2
B3 7 8 jjmit area=B3
IB1 0 4 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
LB1 3 4 LB1
LB2 7 9 LB2
L1 a 1 L1
L2 1 0 L2
L3 1 2 L3
L4 3 5 L4
L5 5 7 L5
L6 7 q L6
LP2 6 0 LP2
LP3 8 0 LP3
RB1 2 102 RB1
LRB1 102 3 LRB1
RB2 5 105 RB2
LRB2 105 0 LRB2
RB3 7 107 RB3
LRB3 107 0 LRB3

.ends



.end


josim -o ./test.csv ./test.cir -V 1
josim-plot.py ./test.csv -t stacked
