master_.param R1   =   5
master_
master_xtest1 one A B Q1
master_xtest2 two Q1 C Q
master_
master_one_.param Lp   =   5
master_one_.param b1   =   1
master_one_.param i1   =   1
master_one_L1 A AA Lp
master_one_L2 B BB 15
master_one_R1 A 0 20
master_one_b1   	30   	10   	 jjmit area=b1
master_one_i1   	0   	30   	pwl(0   	0   	5p   	i1)
master_one_xtest3 three AA BB
master_one_
master_one_three_.param Lp   =   5
master_one_three_.param b1   =   1
master_one_three_.param i1   =   1
master_one_three_L1 25 Ax Lp
master_one_three_L2 15 Bx 15
master_one_three_R1 Bx 0 20
master_one_three_b1   	30   	10   	 jjmit area=b1
master_one_three_i1   	0   	30   	pwl(0   	0   	5p   	i1)
*.ends


two_.param Lp   =   5
two_.param b1   =   1
two_.param i1   =   1
two_L1 0 A Lp
two_L2 15 B 15
two_R1 15 Q 20
two_b1   	30   	10   	 jjmit area=b1
two_i1   	0   	30   	pwl(0   	0   	5p   	i1)
*.ends
