* DSFQ Self clocked Multiplexor
* Author: Adriaan van Wijk
* Version: 1.0
* Last modification date: 21 June 2022
* Last modification by: Adriaan van Wijk
* This testbench uses cells from LS's library of RSFQ cells. This was the version that was tested for layout.

.include cells\LSmitll_DCSFQ_v2p1_optimized.cir
.include cells\LSmitll_JTL_v2p1_optimized.cir
.include AW_TEST_DSFQ_NOT.cir


.param cval=600u

*SO has 10ps of skew here.
I_a0 0 I_a0 pwl(0 0 100p 0 103p cval 105p 0 300p 0 303p cval 305p 0)
I_s0 0 I_s0 pwl(0 0 110p 0 113p cval 115p 0 415p 0 418p cval 420p 0)

.tran 0.25p 500p 0 0.01p

Xsrc_a0 LSmitll_DCSFQ i_a0 src_a0
Xsrc_s0 LSmitll_DCSFQ i_s0 src_s0

Xload_a0 LSMITLL_JTL src_a0 A0
Xload_s0 LSMITLL_JTL src_s0 S0


XNOT DSFQ_NOT A0 S0 Q
* XLOOPA  DSFQ_LOOP   A0      ALOOP
* XLOOPS  DSFQ_LOOP   S0      SLOOP
* XNOT    LSMITLL_NOT ALOOP   SLOOP   Q

Xload_out LSMITLL_JTL Q Qout

Rload Qout 0 2
.print v(A0) v(A1.XNOT) v(A2.XNOT) v(S0) v(CLK2.XNOT) v(Q)

* *$Ports    A B q
* *SFQ PULSE DYNAMIC STORAGE LOOP - Single Time Constant
* .subckt DSFQ_LOOP in q
* .model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)

* *8ps HOLD TIME
* .param LD = 6.5p
* .param RD = 70
* .param RS = 70

* LD in leak LD
* RD leak d1 RD
* RS leak out RS

* BD d1 out jjmit area=0.7
* RBD d1 gg 9.7999
* LBD gg out 5.5369p

* BS leak out jjmit area=1
* RBS leak g9 6.8599
* LBS g9 out 3.8758p
* ROUT out q 0
* .ends


.end