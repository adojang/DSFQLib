* JSIM deck file generated with TimEx
* === DEVICE-UNDER-TEST ===

* === SOURCE DEFINITION ===
.SUBCKT SOURCECELL  8 11
b1   1  2  jjmitll100 area=2.25
b2   3  4  jjmitll100 area=2.25
b3   5  6  jjmitll100 area=2.5
ib1  0  2  pwl(0 0 5p 275ua)
ib2  0  5  pwl(0 0 5p 175ua)
l1   8  7  1p
l2   7  0  3.9p
l3   7  1  0.6p
l4   2  3  1.1p
l5   3  5  4.5p
l6   5  11 2p
lp2  4  0  0.2p
lp3  6  0  0.2p
lrb1 9  2  1p
lrb2 10 4  1p
lrb3 12 6  1p
rb1  1  9  4.31
rb2  3  10 4.31
rb3  5  12 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS SOURCECELL
* === INPUT LOAD DEFINITION ===
.SUBCKT LOADINCELL  2 5
b1 1 6 jjmitll100 area=2.5
b2 4 8 jjmitll100 area=2.5
ib1 0 3 pwl(0 0 5p 350ua)
l1 2 1 2p
l2 1 3 2p
l3 3 4 2p
l4 4 5 2p
lb1 7 6 1p
lb2 9 8 1p
lp1 6 0 0.2p
lp2 8 0 0.2p
rb1 1 7 3.88
rb2 4 9 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS LOADINCELL
* === OUTPUT LOAD DEFINITION ===
.SUBCKT LOADOUTCELL  2 5
b1 1 6 jjmitll100 area=2.5
b2 4 8 jjmitll100 area=2.5
ib1 0 3 pwl(0 0 5p 350ua)
l1 2 1 2p
l2 1 3 2p
l3 3 4 2p
l4 4 5 2p
lb1 7 6 1p
lb2 9 8 1p
lp1 6 0 0.2p
lp2 8 0 0.2p
rb1 1 7 3.88
rb2 4 9 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS LOADOUTCELL
* === SINK DEFINITION ===
.SUBCKT SINKCELL  1
r1 1 0 2
.ENDS SINKCELL
* ===== MAIN ===============================================================================
.param cval=600u

I_gg 0 1000 pwl(0 0 91p 0 94p cval 96p 0)
Rlol 1001 0 2
I_a 0 1001 pwl(0 0 
+100p 0 103p cval 105p 0 
+110p 0 113p cval 115p 0
+300p 0 303p cval 305p 0
+320p 0 323p cval 325p 0
+500p 0 503p cval 505p 0
+530p 0 533p cval 535p 0
+700p 0 703p cval 705p 0
*+740p 0 743p cval 745p 0
+900p 0 903p cval 905p 0
+950p 0 953p cval 955p 0)




XSOURCEINa SOURCECELL 1000 2000
XLOADINa LOADINCELL 2000 A

*XDCSFQ LSmitll_DCSFQ 1000 2000
*XSOURCEINb SOURCECELL 4000 5000
*XLOADINb LOADINCELL 5000 B
XLOADOUTq LOADOUTCELL q xd1
Rcon2 xd1 8000 0
XSINKOUTq SINKCELL 8000



.tran 0.25p 300p 0 0.01p
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)

*$Ports    A B q
*.subckt DSFQ_AND A q
*SFQ PULSE DYNAMIC STORAGE LOOP - Single Time Constant


*Current TAU Try TAU = 10, 20, 30p

*Very sensitive to L1 and RL.
*If BS does not trigger, decrease LD to supply more current to circuit in a shorter timeframe.

* 8 * 0.25 == 2.07ish.
* 0.1 *

*About an 8ps hold time.
*.param LD = 6.5p
*.param RD = 70
*.param RS = 70

*Original Values for atime of about 150ps.
 *.param LD = 5.8p
 .param RD = 6.26
 .param RS = 6.26


.param LD = 7.8p
*.param Rval = 0.4
*.param RD = rval
*.param RS = rval

LD A B LD
RD B C RD
RS B D RS





*The shunted resistor across BD affects the other once since they just combine in paralell. This should be taken into account when doing another review of the NOT gate....



BD C D jjmit area=0.7
RBD C gg 9.7999
LBD gg D 5.5369p


BS B D jjmit area=1
RBS B g9 6.8599
LBS g9 D 3.8758p

*Rcon D q 0

ROUT D q 0

*.print p(A) i(LD) p(B) p(D)

*.print p(A) p(B) p(C) p(D) i(BS) i(RS) i(BD) i(RD) v(B) v(D)
.print i(LD) i(BD) i(BS) i(ROUT) p(BD)

*.print p(A) i(LD) p(B) i(BS) i(BD) i(RS) i(RD) p(D)
*.print i(LD) p(B) i(BS) i(BD) i(RS) i(RD) p(D) i(Rcon)

*.print v(A) i(ROUT) p(A) p(D)

*.print i(LD) i(RD) i(BD) p(D) p(BD) p(BS)
*.print i(LD) i(RD) i(BS) i(RS) p(B) p(D) v(D) i(Rcon)
*.print i(LD) i(BS) i(RD) i(BD) i(RS) p(BS) i(Rcon) v(Rcon)
*.print i(LD) i(RD) i(BS) i(RS) p(B) p(D) p(BD) p(BS)
*.print i(LD) i(RD) i(BS) i(RS)
*.print i(Btest) p(Btest)

*.ends


**************************************** DC TO SFQ **********************************8


* Back-annotated simulation file written by InductEx v.6.0.4 on 2-6-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 2 June 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports 			a q
.subckt LSmitll_DCSFQ a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1.0
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LB=2p
.param LP=0.2p

.param B1=2.25
.param B2=2.25
.param B3=2.5
.param L1=1p
.param L2=3.9p
.param L3=0.6p
.param L4=1.1p
.param L5=4.5p
.param L6=2p
.param IB1=275u
.param IB2=175u
.param LB1=LB
.param LB2=LB
.param LP2=LP
.param LP3=LP
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet

B1 2 3 jjmit area=B1
B2 5 6 jjmit area=B2
B3 7 8 jjmit area=B3
IB1 0 4 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
LB1 3 4 3.12E-12
LB2 7 9 2.281E-12
L1 a 1 1.295E-12
L2 1 0 3.904E-12
L3 1 2 5.998E-13
L4 3 5 1.095E-12
L5 5 7 4.448E-12
L6 7 q 1.334E-12
LP2 6 0 5.16E-13
LP3 8 0 4.733E-13
RB1 2 102 RB1
LRB1 102 3 LRB1
RB2 5 105 RB2
LRB2 105 0 LRB2
RB3 7 107 RB3
LRB3 107 0 LRB3
.ends


.end
