.title KiCad schematic
I2 GND /9 pwl(0 0 5p REF)
L10 /9 /10 Inductor
L9 /5 /9 Inductor
B10 /6 /5 jjmit
LP5 /6 GND Inductor
L8 CLK /5 Inductor
L6 /30 CLK Inductor
B8 /30 /31 jjmit
LP4 /31 GND Inductor
L11 /10 /11 Inductor
B14 /8 /12 jjmit
LP7 /8 GND Inductor
B13 /12 /4 jjmit
I3 GND /4 pwl(0 0 5p REF)
L12 A /4 Inductor
B12 /12 /11 jjmit
LP6 /7 GND Inductor
B11 /7 /10 jjmit
L13 /12 /13 Inductor
L14 /13 /16 Inductor
B16 /15 /17 jjmit
LP9 /15 GND Inductor
LP8 /14 GND Inductor
B15 /14 /13 jjmit
I4 GND /16 pwl(0 0 5p REF)
L15 /16 /17 Inductor
L16 /17 Q Inductor
B9 /24 /23 jjmit
L7 /22 /23 Inductor
L4 /30 /20 Inductor
LP2 /6 GND Inductor
B6 /6 /4 jjmit
B5 /4 /10 jjmit
L3 /10 /30 Inductor
LP3 /24 GND Inductor
B7 /24 /20 jjmit
R2 /22 /20 Resistor
L5 /21 /24 Inductor
R1 /21 /20 Resistor
B3 /3 /10 jjmit
B2 /4 /2 jjmit
L2 B /2 Inductor
B1 /3 /1 jjmit
L1 A /1 Inductor
LP1 /5 GND Inductor
B4 /5 /3 jjmit
I1 GND /10 pwl(0 0 100u)
.end
