.subckt DSFQ_NOT A B C Q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
*A is inverting input.
*B and C are inputs for the OR gate.
*Q is output.

* XDSFQ_OR DSFQ_OR B C CLK
* XJTLCLK LSMITLL_JTLi CLK CLK1
* XNOTLS LSMITLL_NOTi A CLK1 Q


LC_NOT_OR_1 B a_NOT_OR 0
LC_NOT_OR_2 C b_NOT_OR 0
LC_NOT_OR_3 CLK q_NOT_OR 0
*OR GATE
.model jjmit_NOT_OR jj(rtype=1_NOT_OR, vg=2.8mV_NOT_OR, cap=0.07pF_NOT_OR, r0=160_NOT_OR, rn=16_NOT_OR, icrit=0.1mA_NOT_OR)

*Confluence Buffer A
.param l1_NOT_OR = 0.001e-12
.param b1_NOT_OR = 1.44497758
.param b3_NOT_OR = 5.41067564
.param b4_NOT_OR = 7.95470698

* AND GATE LOOP
.param l4_NOT_OR = 1.22182342e-12
.param b7_NOT_OR = 1.59265113
.param b9_NOT_OR = 5.40924075e-01
.param l7_NOT_OR = 1.62539785e-13
.param r1_NOT_OR = 1.09745275e+01
.param r2_NOT_OR = 5.58089917e-01
.param l5_NOT_OR = 5.61756493e-13

* Output Stage
.param b8_NOT_OR = 4.73543077e-01
.param i1_NOT_OR = 3.40214819e-04
.param l3_NOT_OR = 2e-12
.param l6_NOT_OR = 3.06315548e-12

*Confluence Buffer B
.param l2_NOT_OR = l1_NOT_OR
.param b2_NOT_OR = b1_NOT_OR
.param b5_NOT_OR = b3_NOT_OR
.param b6_NOT_OR = b4_NOT_OR

*Parasitics
.param lp1_NOT_OR = 0.2e-12
.param lp2_NOT_OR = 0.2e-12
.param lp3_NOT_OR = 0.2e-12
.param lp4_NOT_OR = 0.2e-12

* Back Annotated .cir file from KiCad
b1_NOT_OR 3_NOT_OR 1_NOT_OR jjmit_NOT_OR area=b1_NOT_OR
b2_NOT_OR 4_NOT_OR 2_NOT_OR jjmit_NOT_OR area=b2_NOT_OR
b3_NOT_OR 3_NOT_OR 10_NOT_OR jjmit_NOT_OR area=b3_NOT_OR
b4_NOT_OR 5_NOT_OR 3_NOT_OR jjmit_NOT_OR area=b4_NOT_OR
b5_NOT_OR 4_NOT_OR 10_NOT_OR jjmit_NOT_OR area=b5_NOT_OR
b6_NOT_OR 6_NOT_OR 4_NOT_OR jjmit_NOT_OR area=b6_NOT_OR
b7_NOT_OR 24_NOT_OR 20_NOT_OR jjmit_NOT_OR area=b7_NOT_OR
b8_NOT_OR 30_NOT_OR 31_NOT_OR jjmit_NOT_OR area=b8_NOT_OR
b9_NOT_OR 24_NOT_OR 23_NOT_OR jjmit_NOT_OR area=b9_NOT_OR
i1_NOT_OR 0 10_NOT_OR pwl(0 0 5p i1_NOT_OR)
l1_NOT_OR a_NOT_OR 1_NOT_OR l1_NOT_OR
l2_NOT_OR b_NOT_OR 2_NOT_OR l2_NOT_OR
l3_NOT_OR 10_NOT_OR 30_NOT_OR l3_NOT_OR
l4_NOT_OR 30_NOT_OR 20_NOT_OR l4_NOT_OR
l5_NOT_OR 21_NOT_OR 24_NOT_OR l5_NOT_OR
l6_NOT_OR 30_NOT_OR q_NOT_OR l6_NOT_OR
l7_NOT_OR 22_NOT_OR 23_NOT_OR l7_NOT_OR
lp1_NOT_OR 5_NOT_OR 0 lp1_NOT_OR
lp2_NOT_OR 6_NOT_OR 0 lp2_NOT_OR
lp3_NOT_OR 24_NOT_OR 0 lp3_NOT_OR
lp4_NOT_OR 31_NOT_OR 0 lp4_NOT_OR
r1_NOT_OR 21_NOT_OR 20_NOT_OR r1_NOT_OR
r2_NOT_OR 22_NOT_OR 20_NOT_OR r2_NOT_OR

*NOT
LC_NOT_NOT_1 A a_NOT1 0
LC_NOT_NOT_2 CLK1 clk_NOT1 0
LC_NOT_NOT_3 Q q_NOT1 0

.model jjmit_NOT1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

.param Phi0_NOT1 = 2.0678e-15
.param B0_NOT1 = 1
.param Ic0_NOT1 = 1.0000e-04
.param IcRs_NOT1 = 6.8599e-04
.param B0Rs_NOT1 = 6.8599
.param Rsheet_NOT1 = 2
.param Lsheet_NOT1 = 1.1300e-12
.param LP_NOT1 = 2.0000e-13
.param IC_NOT1 = 2.5000
.param LB_NOT1 = 2.0000e-12
.param BiasCoef_NOT1 = 0.7000
.param B1_NOT1 = 2.5000
.param B2_NOT1 = 2.5700
.param B3_NOT1 = 1.0700
.param B4_NOT1 = 2.5000
.param B5_NOT1 = 1.3400
.param B6_NOT1 = 3.0300
.param B7_NOT1 = 1.3800
.param B8_NOT1 = 0.8000
.param B9_NOT1 = 2.5000
.param IB1_NOT1 = 1.7500e-04
.param IB2_NOT1 = 8.7000e-05
.param IB3_NOT1 = 2.5700e-04
.param IB4_NOT1 = 1.7500e-04
.param IB5_NOT1 = 1.7500e-04
.param LB1_NOT1 = 2.0000e-12
.param LB2_NOT1 = 2.0000e-12
.param LB3_NOT1 = 2.0000e-12
.param LB4_NOT1 = 2.0000e-12
.param LB5_NOT1 = 2.0000e-12
.param RB1_NOT1 = 2.7440
.param RB2_NOT1 = 2.6692
.param RB3_NOT1 = 6.4111
.param RB4_NOT1 = 2.7440
.param RB5_NOT1 = 5.1193
.param RB6_NOT1 = 2.2640
.param RB7_NOT1 = 4.9709
.param RB8_NOT1 = 8.5749
.param RB9_NOT1 = 2.7440
.param LRB1_NOT1 = 1.5503e-12
.param LRB2_NOT1 = 1.5081e-12
.param LRB3_NOT1 = 3.6223e-12
.param LRB4_NOT1 = 1.5503e-12
.param LRB5_NOT1 = 2.8924e-12
.param LRB6_NOT1 = 1.2792e-12
.param LRB7_NOT1 = 2.8086e-12
.param LRB8_NOT1 = 4.8448e-12
.param LRB9_NOT1 = 1.5503e-12
.param RD_NOT1 = 4
.param LRD_NOT1 = 2.0000e-12

B1_NOT1 1_NOT1 2_NOT1 jjmit_NOT1 area=B1_NOT1
B2_NOT1 4_NOT1 5_NOT1 jjmit_NOT1 area=B2_NOT1
B3_NOT1 7_NOT1 8_NOT1 jjmit_NOT1 area=B3_NOT1
B4_NOT1 13_NOT1 14_NOT1 jjmit_NOT1 area=B4_NOT1
B5_NOT1 17_NOT1 18_NOT1 jjmit_NOT1 area=B5_NOT1
B6_NOT1 10_NOT1 11_NOT1 jjmit_NOT1 area=B6_NOT1
B7_NOT1 20_NOT1 18_NOT1 jjmit_NOT1 area=B7_NOT1
B8_NOT1 18_NOT1 19_NOT1 jjmit_NOT1 area=B8_NOT1
B9_NOT1 21_NOT1 22_NOT1 jjmit_NOT1 area=B9_NOT1

IB1_NOT1 0 3_NOT1 pwl(0 0 5p IB1_NOT1)
IB2_NOT1 0 6_NOT1 pwl(0 0 5p IB2_NOT1)
IB3_NOT1 0 9_NOT1 pwl(0 0 5p IB3_NOT1)
IB4_NOT1 0 15_NOT1 pwl(0 0 5p IB4_NOT1)
IB5_NOT1 0 23_NOT1 pwl(0 0 5p IB5_NOT1)

LB1_NOT1 3_NOT1 1_NOT1 LB1_NOT1
LB2_NOT1 6_NOT1 4_NOT1 LB2_NOT1
LB3_NOT1 8_NOT1 9_NOT1 LB3_NOT1
LB4_NOT1 13_NOT1 15_NOT1 LB4_NOT1
LB5_NOT1 21_NOT1 23_NOT1 LB5_NOT1

L1_NOT1 a_NOT1 1_NOT1 2.062E-12
L2_NOT1 1_NOT1 4_NOT1 1.889E-12
L3_NOT1 4_NOT1 7_NOT1 2.72E-12
L4_NOT1 clk_NOT1 13_NOT1 2.057E-12
L5_NOT1 13_NOT1 16_NOT1 1.029E-12
L6_NOT1 16_NOT1 17_NOT1 1.241E-12
L7_NOT1 16_NOT1 12_NOT1 1.973E-12
L8_NOT1 10_NOT1 12_NOT1 1.003E-12
L9_NOT1 10_NOT1 8_NOT1 7.524E-12
L10_NOT1 8_NOT1 20_NOT1 1.234E-12
L11_NOT1 18_NOT1 21_NOT1 2.607E-12
L12_NOT1 21_NOT1 q_NOT1 2.062E-12

LP1_NOT1 2_NOT1 0 5.271E-13
LP2_NOT1 5_NOT1 0 5.237E-13
LP4_NOT1 14_NOT1 0 4.759E-13
LP6_NOT1 11_NOT1 0 5.021E-13
LP8_NOT1 19_NOT1 0 6.33E-13
LP9_NOT1 22_NOT1 0 4.749E-13

RB1_NOT1 1_NOT1 101_NOT1 RB1_NOT1
LRB1_NOT1 101_NOT1 0 LRB1_NOT1
RB2_NOT1 4_NOT1 104_NOT1 RB2_NOT1
LRB2_NOT1 104_NOT1 5_NOT1 LRB2_NOT1
RB3_NOT1 7_NOT1 107_NOT1 RB3_NOT1
LRB3_NOT1 107_NOT1 8_NOT1 LRB3_NOT1
RB4_NOT1 13_NOT1 113_NOT1 RB4_NOT1
LRB4_NOT1 113_NOT1 0 LRB4_NOT1
RB5_NOT1 17_NOT1 117_NOT1 RB5_NOT1
LRB5_NOT1 117_NOT1 18_NOT1 LRB5_NOT1
RB6_NOT1 10_NOT1 110_NOT1 RB6_NOT1
LRB6_NOT1 110_NOT1 0 LRB6_NOT1
RB7_NOT1 20_NOT1 120_NOT1 RB7_NOT1
LRB7_NOT1 120_NOT1 18_NOT1 LRB7_NOT1
RB8_NOT1 18_NOT1 118_NOT1 RB8_NOT1
LRB8_NOT1 118_NOT1 0 LRB8_NOT1
RB9_NOT1 21_NOT1 121_NOT1 RB9_NOT1
LRB9_NOT1 121_NOT1 0 LRB9_NOT1
LRD_NOT1 12_NOT1 112_NOT1 LRD_NOT1
RD_NOT1 112_NOT1 0 RD_NOT1
* .ends



*JTLNOT
LC_JTLNOT_1 CLK a_JTLNOT 0
LC_JTLNOT_2 CLK1 q_JTLNOT 0

.model jjmit_JTLNOT jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLNOT = 2.0678e-15
.param B0_JTLNOT = 1
.param Ic0_JTLNOT = 1.0000e-04
.param IcRs_JTLNOT = 6.8599e-04
.param B0Rs_JTLNOT = 6.8599
.param Rsheet_JTLNOT = 2
.param Lsheet_JTLNOT = 1.1300e-12
.param LP_JTLNOT = 2.0000e-13
.param IC_JTLNOT = 2.5000
.param Lptl_JTLNOT = 2.0000e-12
.param LB_JTLNOT = 2.0000e-12
.param BiasCoef_JTLNOT = 0.7000
.param B1_JTLNOT = 2.5000
.param B2_JTLNOT = 2.5000
.param IB1_JTLNOT = 3.5000e-04
.param LB1_JTLNOT = 2.0000e-12
.param L1_JTLNOT = 2.0678e-12
.param L2_JTLNOT = 2.0678e-12
.param L3_JTLNOT = 2.0678e-12
.param L4_JTLNOT = 2.0678e-12
.param RB1_JTLNOT = 2.7440
.param RB2_JTLNOT = 2.7440
.param LRB1_JTLNOT = 1.7503e-12
.param LRB2_JTLNOT = 1.7503e-12
.param LP1_JTLNOT = 2.0000e-13
.param LP2_JTLNOT = 2.0000e-13

B1_JTLNOT 1_JTLNOT 2_JTLNOT jjmit_JTLNOT area=B1_JTLNOT
B2_JTLNOT 6_JTLNOT 7_JTLNOT jjmit_JTLNOT area=B2_JTLNOT
IB1_JTLNOT 0 5_JTLNOT pwl(0 0 5p IB1_JTLNOT)
L1_JTLNOT a_JTLNOT 1_JTLNOT 2.082E-12
L2_JTLNOT 1_JTLNOT 4_JTLNOT 2.06E-12
L3_JTLNOT 4_JTLNOT 6_JTLNOT 2.067E-12
L4_JTLNOT 6_JTLNOT q_JTLNOT 2.075E-12
LP1_JTLNOT 2_JTLNOT 0 4.998E-13
LP2_JTLNOT 7_JTLNOT 0 5.011E-13
LB1_JTLNOT 5_JTLNOT 4_JTLNOT LB1_JTLNOT
RB1_JTLNOT 1_JTLNOT 3_JTLNOT RB1_JTLNOT
RB2_JTLNOT 6_JTLNOT 8_JTLNOT RB2_JTLNOT
LRB1_JTLNOT 3_JTLNOT 0 LRB1_JTLNOT
LRB2_JTLNOT 8_JTLNOT 0 LRB2_JTLNOT


.ends
