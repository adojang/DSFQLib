* Author: Adriaan van Wijk
* Version: 1.0
* Last modification date: 21 Feburary 2021
* Last modification by: Adriaan van Wijk

* Copyright (c) 2021 Adriaan van Wijk, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Adriaan van Wijk, 21786275@sun.ac.za


*$Ports 		 A B q
.subckt DSFQ_OR A B q

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

.param Bps=4.50885164e-01
.param Bp=6.38677328e-01
.param Bia=1.08143184e+00
.param Bib=1.20932138e+00
.param Bua=1.03647091e+00
.param Bub=1.10293987e+00
.param Bla=1.56845090e+00
.param Blb= 1.21746914e+00
.param Blim= 1.79155775e+00  
.param LBias =3.15085312e-10
.param Lpoff = 1.30321000e-11
.param Rs=8.18357111e-01
.param RH= 3.64365918e+00
.param IB1= 9.95006250e-05
.param parasitic_induct = 1p

Bia A 1 jjmit area=Bia
Bib B 3 jjmit area=Bib
Bua 1 2 jjmit area=Bua
Bub 3 2 jjmit area=Bub
Bla 1 0 jjmit area=Bla
Blb 3 0 jjmit area=Blb
Bp 4 0 jjmit area=Bp
Bps 5 0 jjmit area=Bps
Blim 6 2 jjmit area=Blim


Ria A 10 1.97
Lia 10 1 parasitic_induct

Rib B 11 1.97
Lib 11 3 parasitic_induct

Rua 1 13 2.16
Lua 13 2 parasitic_induct

Rub 3 14 2.16
Lub 14 2 parasitic_induct

Rla 1 15 1.90
Lla 15 0 parasitic_induct

Rlb 3 16 1.90
Llb 16 0 parasitic_induct

Lpoff 2 4 Lpoff
Rs 4 5 Rs
RH 4 0 RH

Rp 4 17 2.59
Lp 17 0 parasitic_induct

Rps 5 18 2.79
Lps 18 0 parasitic_induct

Lbias VDD 6 Lbias

IB1 0 VDD pwl(0 0 5p IB1 )

Rlim 6 60 1.6
Llim 60 2 parasitic_induct

Lout 2 q 2p
.ends