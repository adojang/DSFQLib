* A Generic Testbench for simulating Logic Gates
* Copyright (c) 2022-2024 Adriaan van Wijk, Stellenbosch University
*
*
* This testbench is not meant to be attached to PTLs as it does not support integrated PTL ports. Basic Circuits Only.


*===== SFQ Source =======
*$Ports 			a q
.subckt LSmitll_DCSFQ a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

.param B0=1.0
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LB=2p
.param LP=0.2p

.param B1=2.25
.param B2=2.25
.param B3=2.5
.param L1=1p
.param L2=3.9p
.param L3=0.6p
.param L4=1.1p
.param L5=4.5p
.param L6=2p
.param IB1=275u
.param IB2=175u
.param LB1=LB
.param LB2=LB
.param LP2=LP
.param LP3=LP
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet

B1 2 3 jjmit area=B1
B2 5 6 jjmit area=B2
B3 7 8 jjmit area=B3
IB1 0 4 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
LB1 3 4 LB1
LB2 7 9 LB2
L1 a 1 L1
L2 1 0 L2
L3 1 2 L3
L4 3 5 L4
L5 5 7 L5
L6 7 q L6
LP2 6 0 LP2
LP3 8 0 LP3
RB1 2 102 RB1
LRB1 102 3 LRB1
RB2 5 105 RB2
LRB2 105 0 LRB2
RB3 7 107 RB3
LRB3 107 0 LRB3

.ends

*=========== JTL LOADS ==========
*$Ports 			a q
.subckt LSMITLL_JTL a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=IC
.param IB1=(B1+B2)*Ic0*BiasCoef
.param LB1=LB
.param L1=Phi0/(4*B1*Ic0)
.param L2=Phi0/(4*B1*Ic0)
.param L3=Phi0/(4*B1*Ic0)
.param L4=Phi0/(4*B2*Ic0)
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP

B1 1 2 jjmit area=B1
B2 6 7 jjmit area=B2
IB1 0 5 pwl(0 0 5p IB1)
L1 a 1 L1
L2 1 4 L2
L3 4 6 L3
L4 6 q L4
LP1 2 0 LP1
LP2 7 0 LP2
LB1 5 4 LB1
RB1 1 3 RB1
RB2 6 8 RB2
LRB1 3 0 LRB1
LRB2 8 0 LRB2

.ends

*====== Device Under Test ======
*$Ports     A B Q
.subckt DUT A B Q

*there should be a dc bias in here somewhere.

.model 50 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=50uA)
.model 70 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=70uA)
.model 100 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)
.model 120 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=120uA)
.model 130 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=130uA)
.model 180 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=180uA)

*Ibias vdd 0 dc 180u

Bia A 1 120
Bib B 3 120

Bua 1 2 100
Bub 3 2 100

Bla 1 0 130
Blb 3 0 130

Lpoff 2 4 16p

Rs 4 5 1

Bp 4 0 70
Bps 5 0 50

Lbias Q 0 350p
Blim 2 Q 180

.ends

*=========== END DUT =========

*====== Main TestBench========


XSourceA LSmitll_DCSFQ srcAin srcAout
XSourceB LSmitll_DCSFQ srcBin srcBout

XLoadInA LSMITLL_JTL srcAout loadaout
XLoadInB LSMITLL_JTL srcBout loadbout

*=======================================
XDUT DUT loadaout loadbout dutout
*=======================================

XLoadCircuit LSMITLL_JTL dutout loadout
RSink loadout 0 2

* ==SOURCE CURRENT INPUTS==

* The tests below are preconfigured for common logic gate tests.
* The tests include timing tests which are neccesary for DSFQ to be verified.
* If two inputs arrive within X time of one another, both are considered (nominally 40ps)

*700u is a good avg value i guess
.param cval = 700u


* BASIC Timing Tests are each 100ps apart:
IsrcA 0 srcAin pwl(0 0 100p 0 101p cval 102p 0 300p 0 201p cval 202p 0)
IsrcB 0 srcBin pwl(0 0 200p 0 201p cval 202p 0 300p 0 201p cval 202p 0)

* BASIC Timing Tests each 50ps apart:
*IsrcA 0 srcAin pwl(0 0 50p 0 51p cval 52p 0 150p 0 151p cval 152p 0)
*IsrcB 0 srcBin pwl(0 0 100p 0 101p cval 102p 0 150p 0 151p cval 152p 0)

* Advanced Tests to see how long a value is held 30ps 40ps 50ps
*IsrcA 0 srcAin pwl(0 0 50p 0 51p cval 52p 0 200p 0 201p cval 202p 0 300p 0 301p cval 302p 0)
*IsrcB 0 srcBin pwl(0 0 80p 0 81p cval 82p 0 240p 0 241p cval 242p 0 350p 0 351p cval 352p 0)


* Advanced Tests to demonstrate multiple input rejection
.tran 0.25p 500p 0 0.25p

*Prints Circuit Inputs, and Circuit Output


.print i(Lpoff.XDUT) i(Lbias.XDUT) p(Bia.XDUT) p(Bib.XDUT) i(Rs.XDUT) p(Blim.XDUT) i(L1.XLoadCircuit) p(B1.XLoadCircuit) i(RSink)
*.print i(L4.XLoadInA) i(L4.XLoadInB)
*.print i(L1.XSourceA) i(L1.XSourceB) i(L6.XSourceA) i(L6.XSourceB)

*Check Sources
*.print i(L6.XSourceA) i(L6.XSourceB) i(L4.XLoadInA) i(L4.XLoadInB)

*Default Input Output Prints
*.print i(L6.XSourceA) i(L6.XSourceB) i(RSink) p(Blim.XDUT) p(B1.XLoadCircuit)

.end