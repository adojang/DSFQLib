.subckt master A B C Q
.PARAM LAD  	=	 	    5

xtest1 one A B Q1
xtest2 two Q1 C Q


.subckt one Am Bm Q1m
L1 Am Bm 5
R1 Am 0 5
C1 Am Qm1

xtest3 three AA BB

.subckt three AA BB
L1 AA BB 55
.ends

.ends


.subckt two Q1m Cm Q
L1 Q1m Cm 5
R1 Q1 0 5
C1 Q11 Q
.ends





.ends