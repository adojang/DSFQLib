* Adapted from DSFQ_AND Gate by Rylov
* Author: AJ. van Wijk
* Version: 1.0
* Last modification date: 25 April 2022
* Last modification by: AJ. van Wijk

.param cval=600u

I_a 0 1000 pwl(0 0 
+100p 0 103p cval 105p 0
+300p 0 303p cval 305p 0
+350p 0 353p cval 355p 0
+400p 0 403p cval 405p 0
+450p 0 453p cval 455p 0
+500p 0 503p cval 505p 0
+710p 0 713p cval 715p 0
+820p 0 823p cval 825p 0
+850p 0 853p cval 855p 0)

I_b 0 4000 pwl(0 0 
+200p 0 203p cval 205p 0
+300p 0 303p cval 305p 0
+350p 0 353p cval 355p 0
+405p 0 408p cval 410p 0
+460p 0 463p cval 465p 0
+515p 0 518p cval 520p 0
+710p 0 713p cval 715p 0
+820p 0 823p cval 825p 0
+850p 0 853p cval 855p 0)

XSOURCEINa LSmitll_DCSFQ 1000 2000
XLOADINa LSMITLL_JTL 2000 A
XSOURCEINb LSmitll_DCSFQ 4000 5000
XLOADINb LSMITLL_JTL 5000 B
XLOADOUTq LSMITLL_JTL q 8000
XLOADDC   LSmitll_SFQDC 8000 9000

Rout 9000 0 2

XDUT DSFQ_AND A B q

.tran 0.25p 600p 0 0.01p
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)

.print v(L1.XLOADINa) v(L1.XLOADINb) v(Rout) p(B5.XDUT)


.subckt DSFQ_AND A B q
*Tuned Parameters
.param l1       =                3.09037291e-12
.param l3       =                2.03058886e-12
.param r1       =                7.04349127e-01
.param r3       =                1.34323634e+00
.param rbias    =                1.00298596e+02

.param l2       =         l1
.param r2       =         r1
.param r4       =         r3

*Static Parameters
.param b1       =         5.16417451e-01
.param b2       =         b1
.param b3       =         3.5e-01
.param b4       =         b3
.param b5       =         1.05188201e+00

.param rb1      =         12.92859137e+00
.param rb2      =         12.92013085e+00
.param rb3      =         19.98871344e+00
.param rb4      =         19.98963516e+00
.param rb5      =         6.566007373e+00

.param lrb1     =         3.94321337e-13
.param lrb2     =         5.33421859e-13
.param lrb3     =         1.39314087e-12
.param lrb4     =         1.41001012e-12
.param lrb5     =         1.19776828e-12
.param lp1      =         8.25215763e-13

b1   	4   	5   	 jjmit area=b1
b2   	6   	7   	 jjmit area=b2
b3   	4   	8   	 jjmit area=b3
b4   	6   	4   	 jjmit area=b4
b5   	4   	9   	 jjmit area=b5
v1   	0   	bias   	pwl(0   	0   	5p   	2.067m)
Rbias   bias    bias1   Rbias
Lbias   bias1   4       12p

l1   	a   	5   	 l1
l2   	b   	7   	 l2
l3   	4   	q   	 l3
lp1   	9   	0   	 lp1
lrb1   	10   	4   	 lrb1
lrb2   	11   	6   	 lrb2
lrb3   	12   	4   	 lrb3
lrb4   	13   	6   	 lrb4
lrb5   	14   	0   	 lrb5
r1   	5   	4   	 r1
r2   	7   	6   	 r2
r3   	8   	5   	 r3
r4   	4   	7   	 r4
rb1   	5   	10   	 rb1
rb2   	7   	11   	 rb2
rb3   	8   	12   	 rb3
rb4   	4   	13   	 rb4
rb5   	4   	14   	 rb5

.ends

.subckt LSMITLL_JTL a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=IC
.param IB1=(B1+B2)*Ic0*BiasCoef
.param LB1=LB
.param L1=Phi0/(4*B1*Ic0)
.param L2=Phi0/(4*B1*Ic0)
.param L3=Phi0/(4*B1*Ic0)
.param L4=Phi0/(4*B2*Ic0)
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP

B1 1 2 jjmit area=B1
B2 6 7 jjmit area=B2
IB1 0 5 pwl(0 0 5p IB1)
L1 a 1 2.082E-12
L2 1 4 2.06E-12
L3 4 6 2.067E-12
L4 6 q 2.075E-12
LP1 2 0 4.998E-13
LP2 7 0 5.011E-13
LB1 5 4 LB1
RB1 1 3 RB1
RB2 6 8 RB2
LRB1 3 0 LRB1
LRB2 8 0 LRB2
.ends


*$Ports 			a q
.subckt LSmitll_DCSFQ a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1.0
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LB=2p
.param LP=0.2p

.param B1=2.25
.param B2=2.25
.param B3=2.5
.param L1=1p
.param L2=3.9p
.param L3=0.6p
.param L4=1.1p
.param L5=4.5p
.param L6=2p
.param IB1=275u
.param IB2=175u
.param LB1=LB
.param LB2=LB
.param LP2=LP
.param LP3=LP
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet

B1 2 3 jjmit area=B1
B2 5 6 jjmit area=B2
B3 7 8 jjmit area=B3
IB1 0 4 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
LB1 3 4 3.12E-12
LB2 7 9 2.281E-12
L1 a 1 1.295E-12
L2 1 0 3.904E-12
L3 1 2 5.998E-13
L4 3 5 1.095E-12
L5 5 7 4.448E-12
L6 7 q 1.334E-12
LP2 6 0 5.16E-13
LP3 8 0 4.733E-13
RB1 2 102 RB1
LRB1 102 3 LRB1
RB2 5 105 RB2
LRB2 105 0 LRB2
RB3 7 107 RB3
LRB3 107 0 LRB3
.ends


*$Ports a q
.subckt LSmitll_SFQDC a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12
.param LB=2p
.param LP=0.5p

.param B1=3.25
.param B2=2.00
.param B3=1.50
.param B4=3.00
.param B5=1.75
.param B6=1.50
.param B7=1.50
.param B8=2.00

.param IB1=280u
.param IB2=150u
.param IB3=220u
.param IB4=80u

.param L1=1.522p
.param L3=0.827p
.param L4=1.12884p
.param L5=1.11098p
.param L5b=3.216p
.param L6=5.94p
.param L10=0.215p
.param L19=0.954p
.param L13=3.699p
.param L18=2.010p
.param L17=1.510p
.param LR1=0.91p
.param R1=0.375

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8

.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LP1=LP
.param LP4=LP
.param LP5=LP
.param LP7=LP
.param LP8=LP

B1 2 4 jjmit area=B1
B2 7 10 jjmit area=B2
B3 6 8 jjmit area=B3
B4 10 11 jjmit area=B4
B5 8 15 jjmit area=B5
B6 17 18 jjmit area=B6
B7 20 21 jjmit area=B7
B8 24 25 jjmit area=B8

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
IB3 0 19 pwl(0 0 5p IB3)
IB4 0 23 pwl(0 0 5p IB4)

LB1 2 3 LB1
LB2 8 9 LB2
LB3 18 19 LB3
LB4 22 23 LB4

L1 a 2 1.402E-12
L3 2 5 8.739E-13
L4 5 6 1.294E-12
L5 5 7 1.307E-12
L5B 10 12 3.216E-12
L6 8 12 5.963E-12
L10 12 17 4.424E-13
L13 20 22 3.547E-12
L17 24 q 1.22E-12
L18 22 24 2.081E-12
L19 18 20 7.952E-13

LR1 12 13 9.02E-13
R1 13 0 R1

LP1 4 0 3.705E-13
LP4 11 0 4.154E-13
LP5 15 0 4.837E-13
LP7 21 0 5.043E-13
LP8 25 0 4.001E-13

RB1 2 102 RB1
LRB1 102 0 LRB1
RB2 7 107 RB2
LRB2 107 10 LRB2
RB3 6 106 RB3
LRB3 106 8 LRB3
RB4 10 110 RB4
LRB4 110 0 LRB4
RB5 8 108 RB5
LRB5 108 0 LRB5
RB6 17 117 RB6
LRB6 117 18 LRB6
RB7 20 120 RB7
LRB7 120 0 LRB7
RB8 24 124 RB8
LRB8 124 0 LRB8
.ends


.end