.title KiCad schematic
LRB5 Net-_LRB5-Pad1_ GND Inductor
LP1 Net-_B5-Pad1_ GND Inductor
LRB4 Net-_LRB4-Pad1_ Net-_B1-Pad1_ Inductor
RB4 Net-_B4-Pad2_ Net-_LRB4-Pad1_ Resistor
RB3 Net-_B3-Pad2_ Net-_LRB3-Pad1_ Resistor
LRB3 Net-_LRB3-Pad1_ Net-_B1-Pad1_ Inductor
RB5 Net-_B1-Pad1_ Net-_LRB5-Pad1_ Resistor
L3 Net-_B1-Pad1_ Q Inductor
B5 Net-_B5-Pad1_ Net-_B1-Pad1_ jjmit
I1 GND Net-_B1-Pad1_ pwl(0 0 5p REF)
L2 B Net-_B2-Pad2_ Inductor
L1 A Net-_B1-Pad2_ Inductor
R3 Net-_B3-Pad2_ Net-_B1-Pad2_ Resistor
RB2 Net-_B2-Pad2_ Net-_LRB2-Pad1_ Resistor
LRB2 Net-_LRB2-Pad1_ Net-_B1-Pad1_ Inductor
B4 Net-_B1-Pad1_ Net-_B4-Pad2_ jjmit
R4 Net-_B4-Pad2_ Net-_B2-Pad2_ Resistor
RB1 Net-_B1-Pad2_ Net-_LRB1-Pad1_ Resistor
LRB1 Net-_LRB1-Pad1_ Net-_B1-Pad1_ Inductor
B3 Net-_B1-Pad1_ Net-_B3-Pad2_ jjmit
R2 Net-_B2-Pad2_ Net-_B1-Pad1_ Resistor
B2 Net-_B1-Pad1_ Net-_B2-Pad2_ jjmit
B1 Net-_B1-Pad1_ Net-_B1-Pad2_ jjmit
R1 Net-_B1-Pad2_ Net-_B1-Pad1_ Resistor
.end
