#Original Parameters for 10ps skew

.param 	b1  	= 0.84
.param 	b2  	= 0.84
.param 	b3  	= 0.6
.param 	b4  	= 0.6
.param 	b5  	= 1.68
.param 	i1  	= 70u
.param 	l1  	= 8p
.param 	l2  	= 8p
.param 	l3  	= 2p
.param 	lp1  	= 0.2p
.param 	lrb1  	= 6.4597p
.param 	lrb2  	= 4.6141p
.param 	lrb3  	= 6.4597p
.param 	lrb4  	= 4.6141p
.param 	lrb5  	= 2.3071p

.param  Rhold   = 3.3248

.param 	rA  	= Rhold
*.param 	r2  	= Rhold
*.param 	r3  	= Rhold
*.param 	r4  	= Rhold

.param 	rb1  	= 11.4332
.param 	rb2  	= 8.1666
.param 	rb3  	= 11.4332
.param 	rb4  	= 8.1666
.param 	rb5  	= 4.0833