.param 	b1  	= 
.param 	b2  	= 
.param 	b3  	= 
.param 	b4  	= 
.param 	b5  	= 
.param 	i1  	= 
.param 	l1  	= 
.param 	l2  	= 
.param 	l3  	= 
.param 	lp1  	= 
.param 	lrb1  	= 
.param 	lrb2  	= 
.param 	lrb3  	= 
.param 	lrb4  	= 
.param 	lrb5  	= 
.param 	r1  	= 
.param 	r2  	= 
.param 	r3  	= 
.param 	r4  	= 
.param 	rb1  	= 
.param 	rb2  	= 
.param 	rb3  	= 
.param 	rb4  	= 
.param 	rb5  	= 


* Back Annotated .cir file from KiCad
b1   	3   	2   	 jjmit area=b1
b2   	3   	4   	 jjmit area=b2
b3   	3   	5   	 jjmit area=b3
b4   	3   	6   	 jjmit area=b4
b5   	7   	3   	 jjmit area=b5
i1   	0   	3   	pwl(0   	0   	5p   	i1)
l1   	a   	2   	 l1
l2   	b   	4   	 l2
l3   	3   	q   	 l3
lp1   	7   	0   	 lp1
lrb1   	8   	3   	 lrb1
lrb2   	9   	3   	 lrb2
lrb3   	10   	3   	 lrb3
lrb4   	11   	3   	 lrb4
lrb5   	12   	0   	 lrb5
r1   	5   	2   	 r1
r2   	6   	4   	 r2
r3   	2   	3   	 r3
r4   	4   	3   	 r4
rb1   	2   	8   	 rb1
rb2   	4   	9   	 rb2
rb3   	5   	10   	 rb3
rb4   	6   	11   	 rb4
rb5   	3   	12   	 rb5
.end