* Author: Adriaan van Wijk
* Version: 1.0
* Last modification date: 21 Feburary 2021
* Last modification by: Adriaan van Wijk
* Based on the design by Rylov [2019]

* Copyright (c) 2021 Adriaan van Wijk, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Adriaan van Wijk, 21786275@sun.ac.za



*$Ports    A B q
.subckt DSFQ_AND A B q
.param pInduc = 1p

.param main=0.84
.param secondary=0.60
.param third=1.68
.param pInduc = 1p
.param retentionResistor=4


.param Ibiasz=70u
.param L1=12p
.param L2=12p 
.param Lout=2p
.param retentionResistor=4


L1 A 1 L1
L2 B 4 L2
RD1 1 2 0.67
RD2 4 5 0.67
BD1 2 C jjmit area=secondary
RDp1 2 14 2.8
Ld1 14 C pInduc
BD2 5 C jjmit area=secondary
RDp2 5 15 2.8
Ld2 15 C pInduc
Rh1 1 C retentionResistor
Rh2 4 C retentionResistor
B1 1 C jjmit area=main
Rb1 1 10 2.37
Lb1 10 C pInduc
B2 4 C jjmit area=main
Rb2 4 11 2.37
Lb2 11 C pInduc
B3 C 0 jjmit area=third
Rb3 C 13 1.67
Lb3 13 0 pInduc
Ibias 0 C dc Ibiasz
Lout C q Lout
.ends