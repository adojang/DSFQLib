.subckt DSFQ_MUX D0 D1 S Q

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=100uA)


* XSPLITA LSMITLL_SPLIT D0 A1 CLK1
* XSPLITS LSMITLL_SPLIT S S1 S3


XJTLA1 LSMITLL_JTL D0 A2a
XJTLA2 LSMITLL_JTL A2a A2


XJTLCLK LSMITLL_JTL D0 CLK1
XJTLCLK2 LSMITLL_JTL CLK1 CLK2




XJTLS1 LSMITLL_JTL S S1
XJTLS3 LSMITLL_JTL S 2
* XJTLS3a LSMITLL_JTL S4a S4

* XJTLB LSMITLL_JTL D1 B1a
XJTLBa LSMITLL_JTL D1 B1

XJTLQ1 LSMITLL_JTL Q1a Q1
XJTLQ2a LSMITLL_JTL Q2a Q2b
XJTLQ2b LSMITLL_JTL Q2b Q2

XAND1   DSFQ_AND   A2 A3 Q1a
XAND2   DSFQ_AND   S2 B1 Q2a
XNOT    DSFQ_NOT S1 CLK2 CLK2 A3
XOR     DSFQ_OR    Q1 Q2 Q


* I_s0 0 Q2a pwl(0 0 5p 100u)
* B_xA1   Q2a   	Q2   	 jjmit area=1.5

* I_s02 0 B1a pwl(0 0 5p 200u)
* B_xA12   B1a   	B1   	 jjmit area=2.5



.ends