.param 	b1  	= 
.param 	b2  	= 
.param 	b3  	= 
.param 	b4  	= 
.param 	b5  	= 
.param 	b6  	= 
.param 	b7  	= 
.param 	b8  	= 
.param 	b9  	= 
.param 	i1  	= 
.param 	l1  	= 
.param 	l2  	= 
.param 	l3  	= 
.param 	l4  	= 
.param 	l5  	= 
.param 	l6  	= 
.param 	l7  	= 
.param 	lp1  	= 
.param 	lp2  	= 
.param 	lp3  	= 
.param 	lp4  	= 
.param 	r1  	= 
.param 	r2  	= 


* Back Annotated .cir file from KiCad
b1   	3   	1   	 jjmit area=b1
b2   	4   	2   	 jjmit area=b2
b3   	3   	10   	 jjmit area=b3
b4   	5   	3   	 jjmit area=b4
b5   	4   	10   	 jjmit area=b5
b6   	6   	4   	 jjmit area=b6
b7   	24   	20   	 jjmit area=b7
b8   	30   	31   	 jjmit area=b8
b9   	24   	23   	 jjmit area=b9
i1   	0   	10   	pwl(0   	0   	100u) i1
l1   	a   	1   	 l1
l2   	b   	2   	 l2
l3   	10   	30   	 l3
l4   	30   	20   	 l4
l5   	21   	24   	 l5
l6   	30   	q   	 l6
l7   	22   	23   	 l7
lp1   	5   	0   	 lp1
lp2   	6   	0   	 lp2
lp3   	24   	0   	 lp3
lp4   	31   	0   	 lp4
r1   	21   	20   	 r1
r2   	22   	20   	 r2
.end