.subckt RYLOV a b q
.param 	b1  	= 0.84
.param 	b2  	= 0.84
.param 	b3  	= 0.60
.param 	b4  	= 0.60
.param 	b5  	= 1.68
.param 	i1  	= 70u
.param 	l1  	= 7p
.param 	l2  	= 7p
.param 	l3  	= 2p
.param 	lp1  	= 0.2p
.param 	lrb5  	= 2.3071p
.param 	r1  	= 4
.param 	r2  	= 4
.param 	r3  	= 0.68
.param 	r4  	= 0.68
.param 	rb5  	= 4.0833

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
* Back Annotated .cir file from KiCad
b1   	10   	39   	 jjmit area=b1
b2   	30   	20   	 jjmit area=b2
b3   	12   	39   	 jjmit area=b3
b4   	30   	22   	 jjmit area=b4
b5   	30m   	31   	 jjmit area=b5
i1   	0   	30m   	pwl(0   	0   	5p   	i1)
l1   	a   	10   	 l1
l2   	b   	20   	 l2
l3   	30m   	q   	 l3
lp1   	31   	0   	 lp1
lrb5   	32   	0   	 lrb5
r1   	10   	39   	 r1

lmeasure      39      30      0
lmeasure2       30      30m   0
r2   	20   	30   	 r2
r3   	12   	10   	 r3
r4   	22   	20   	 r4
rb5   	30m   	32   	 rb5
.ends