* Author: A. van Wijk
* Version: 1.0
* Last modification date: 09 January 2023
* Last modification by: A. van Wijk
* Copyright (c) 2022 Adriaan van Wijk, Stellenbosch University
* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:
* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.
* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Adriaan van Wijk, jacowijka@gmail.com
* The cell is not designed to be connected directly to passive transmission lines
* The cell is designed for a skew time of 8ps. 
* Maximum system clock speed of 125GHz

.subckt DSFQ_ANDx a b q
.param 	b1  	= 0.84
.param 	b2  	= 0.84
.param 	b3  	= 0.60
.param 	b4  	= 0.60
.param 	b5  	= 1.68
.param 	i1  	= 70u
.param 	l1  	= 2p
.param 	l2  	= 4p
.param 	l3  	= 2p
.param 	lp1  	= 0.2p
.param 	lrb5  	= 2.3071p
.param 	r1  	= 4
.param 	r2  	= 4
.param 	r3  	= 0.68
.param 	r4  	= 0.68
.param 	rb5  	= 4.0833

.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
* Back Annotated .cir file from KiCad
b1   	10   	30   	 jjmit area=b1
b2   	30   	20   	 jjmit area=b2
b3   	12   	30   	 jjmit area=b3
b4   	30   	22   	 jjmit area=b4
b5   	30   	31   	 jjmit area=b5
i1   	0   	30   	pwl(0   	0   	5p   	i1)
l1   	a   	10   	 l1
l2   	b   	20   	 l2
l3   	30   	q   	 l3
lp1   	31   	0   	 lp1
lrb5   	32   	0   	 lrb5
r1   	10   	30   	 r1



r2   	20   	30   	 r2
r3   	12   	10   	 r3
r4   	22   	20   	 r4
rb5   	30   	32   	 rb5
.ends