.param 	b1  	= 1.2
.param 	b2  	= 1.2
.param 	b3  	= 1
.param 	b4  	= 1.3
.param 	b5  	= 1
.param 	b6  	= 1.3
.param 	b7  	= 0.7
.param 	b8  	= 1.8
.param 	b9  	= 0.5
.param 	i1  	= 250u
.param 	l1  	= 2p
.param 	l2  	= 2p
.param 	l3  	= 4p
.param 	l4  	= 16p
.param 	l5  	= 350p
.param 	lp4  	= 1p
.param 	lp6  	= 1p
.param 	lp7  	= 1p
.param 	lp9  	= 1p
.param 	lrb1  	= 3.229p
.param 	lrb2  	= lrb1
.param 	lrb3  	= 3.8758p
.param 	lrb4  	= 2.9814p
.param 	lrb5  	= lrb3
.param 	lrb6  	= lrb4
.param 	lrb7  	= 5.5369p
.param 	lrb8  	= 2.1532p
.param 	lrb9  	= 7.7517p
.param 	r1  	= 1
.param 	rb1  	= 5.7166
.param 	rb2  	= rb1
.param 	rb3  	= 6.8599
.param 	rb4  	= 5.2768
.param 	rb5  	= rb3
.param 	rb6  	= rb4
.param 	rb7  	= 9.799
.param 	rb8  	= 3.811
.param 	rb9  	= 13.7198


* Back Annotated .cir file from KiCad
b1   	2   	3   	 jjmit area=b1
b2   	4   	5   	 jjmit area=b2
b3   	2   	6   	 jjmit area=b3
b4   	7   	2   	 jjmit area=b4
b5   	4   	6   	 jjmit area=b5
b6   	8   	4   	 jjmit area=b6
b7   	9   	10   	 jjmit area=b7
b8   	11   	q   	 jjmit area=b8
b9   	12   	13   	 jjmit area=b9
i1   	0   	6   	pwl(0   	0   	100u) i1
l1   	a   	3   	 l1
l2   	b   	5   	 l2
l3   	6   	q   	 l3
l4   	q   	10   	 l4
l5   	11   	0   	 l5
lp4   	7   	0   	 lp4
lp6   	8   	0   	 lp6
lp7   	9   	0   	 lp7
lp9   	12   	0   	 lp9
lrb1   	14   	2   	 lrb1
lrb2   	15   	4   	 lrb2
lrb3   	16   	2   	 lrb3
lrb4   	17   	0   	 lrb4
lrb5   	18   	4   	 lrb5
lrb6   	19   	0   	 lrb6
lrb7   	20   	0   	 lrb7
lrb8   	21   	11   	 lrb8
lrb9   	22   	0   	 lrb9
r1   	10   	13   	 r1
rb1   	3   	14   	 rb1
rb2   	5   	15   	 rb2
rb3   	6   	16   	 rb3
rb4   	2   	17   	 rb4
rb5   	6   	18   	 rb5
rb6   	4   	19   	 rb6
rb7   	10   	20   	 rb7
rb8   	q   	21   	 rb8
rb9   	13   	22   	 rb9
.end