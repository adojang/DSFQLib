*This Subcircuit was flattened. The AND gate has a slightly smaller output inductance than is typical, which may change the normal margins.


.subckt DSFQ_XOR A B Q

* XSPLITA LSmitll_SPLITo A A1 A2
* XSPLITB LSmitll_SPLITo B B1 B2

* XJTL1 LSmitll_JTLi A1 A11
* XJTL2 LSmitll_JTLi B1 B11
* XJTL3 LSmitll_JTLi OR1 OR2
* XJTL4 LSmitll_JTLi OR2 OR3

* XNAND1  DSFQ_ANDo    A1     B1   AND1
* XNAND2  DSFQ_NOTo    AND1   A11   B11   AND2
* XOR     DSFQ_ORi     A1     B2   OR1
* XAND    DSFQ_ANDo    AND2   OR3  Q

*Libraries so the circuit can run by itself without requiring the user to add them.
*Libraries Included: DSFQ_AND DSFQ_OR LSMITLL_JTL, LSMITLL_SPLIT, LSMITLL_NOT DSFQ_NOT, 


*****JTL CELLS ***********************************************
*JTLA1
LC_JTLA1_1 A1 a_JTLA1 0
LC_JTLA1_2 A11 q_JTLA1 0

.model jjmit_JTLA1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLA1 = 2.0678e-15
.param B0_JTLA1 = 1
.param Ic0_JTLA1 = 1.0000e-04
.param IcRs_JTLA1 = 6.8599e-04
.param B0Rs_JTLA1 = 6.8599
.param Rsheet_JTLA1 = 2
.param Lsheet_JTLA1 = 1.1300e-12
.param LP_JTLA1 = 2.0000e-13
.param IC_JTLA1 = 2.5000
.param Lptl_JTLA1 = 2.0000e-12
.param LB_JTLA1 = 2.0000e-12
.param BiasCoef_JTLA1 = 0.7000
.param B1_JTLA1 = 2.5000
.param B2_JTLA1 = 2.5000
.param IB1_JTLA1 = 3.5000e-04
.param LB1_JTLA1 = 2.0000e-12
.param L1_JTLA1 = 2.0678e-12
.param L2_JTLA1 = 2.0678e-12
.param L3_JTLA1 = 2.0678e-12
.param L4_JTLA1 = 2.0678e-12
.param RB1_JTLA1 = 2.7440
.param RB2_JTLA1 = 2.7440
.param LRB1_JTLA1 = 1.7503e-12
.param LRB2_JTLA1 = 1.7503e-12
.param LP1_JTLA1 = 2.0000e-13
.param LP2_JTLA1 = 2.0000e-13

B1_JTLA1 1_JTLA1 2_JTLA1 jjmit_JTLA1 area=B1_JTLA1
B2_JTLA1 6_JTLA1 7_JTLA1 jjmit_JTLA1 area=B2_JTLA1
IB1_JTLA1 0 5_JTLA1 pwl(0 0 5p IB1_JTLA1)
L1_JTLA1 a_JTLA1 1_JTLA1 2.082E-12
L2_JTLA1 1_JTLA1 4_JTLA1 2.06E-12
L3_JTLA1 4_JTLA1 6_JTLA1 2.067E-12
L4_JTLA1 6_JTLA1 q_JTLA1 2.075E-12
LP1_JTLA1 2_JTLA1 0 4.998E-13
LP2_JTLA1 7_JTLA1 0 5.011E-13
LB1_JTLA1 5_JTLA1 4_JTLA1 LB1_JTLA1
RB1_JTLA1 1_JTLA1 3_JTLA1 RB1_JTLA1
RB2_JTLA1 6_JTLA1 8_JTLA1 RB2_JTLA1
LRB1_JTLA1 3_JTLA1 0 LRB1_JTLA1
LRB2_JTLA1 8_JTLA1 0 LRB2_JTLA1

*JTLA2
LC_JTLA2_1 B1 a_JTLA2 0
LC_JTLA2_2 B11 q_JTLA2 0

.model jjmit_JTLA2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLA2 = 2.0678e-15
.param B0_JTLA2 = 1
.param Ic0_JTLA2 = 1.0000e-04
.param IcRs_JTLA2 = 6.8599e-04
.param B0Rs_JTLA2 = 6.8599
.param Rsheet_JTLA2 = 2
.param Lsheet_JTLA2 = 1.1300e-12
.param LP_JTLA2 = 2.0000e-13
.param IC_JTLA2 = 2.5000
.param Lptl_JTLA2 = 2.0000e-12
.param LB_JTLA2 = 2.0000e-12
.param BiasCoef_JTLA2 = 0.7000
.param B1_JTLA2 = 2.5000
.param B2_JTLA2 = 2.5000
.param IB1_JTLA2 = 3.5000e-04
.param LB1_JTLA2 = 2.0000e-12
.param L1_JTLA2 = 2.0678e-12
.param L2_JTLA2 = 2.0678e-12
.param L3_JTLA2 = 2.0678e-12
.param L4_JTLA2 = 2.0678e-12
.param RB1_JTLA2 = 2.7440
.param RB2_JTLA2 = 2.7440
.param LRB1_JTLA2 = 1.7503e-12
.param LRB2_JTLA2 = 1.7503e-12
.param LP1_JTLA2 = 2.0000e-13
.param LP2_JTLA2 = 2.0000e-13

B1_JTLA2 1_JTLA2 2_JTLA2 jjmit_JTLA2 area=B1_JTLA2
B2_JTLA2 6_JTLA2 7_JTLA2 jjmit_JTLA2 area=B2_JTLA2
IB1_JTLA2 0 5_JTLA2 pwl(0 0 5p IB1_JTLA2)
L1_JTLA2 a_JTLA2 1_JTLA2 2.082E-12
L2_JTLA2 1_JTLA2 4_JTLA2 2.06E-12
L3_JTLA2 4_JTLA2 6_JTLA2 2.067E-12
L4_JTLA2 6_JTLA2 q_JTLA2 2.075E-12
LP1_JTLA2 2_JTLA2 0 4.998E-13
LP2_JTLA2 7_JTLA2 0 5.011E-13
LB1_JTLA2 5_JTLA2 4_JTLA2 LB1_JTLA2
RB1_JTLA2 1_JTLA2 3_JTLA2 RB1_JTLA2
RB2_JTLA2 6_JTLA2 8_JTLA2 RB2_JTLA2
LRB1_JTLA2 3_JTLA2 0 LRB1_JTLA2
LRB2_JTLA2 8_JTLA2 0 LRB2_JTLA2

*JTLA3
LC_JTLA3_1 OR1 a_JTLA3 0
LC_JTLA3_2 OR2 q_JTLA3 0

.model jjmit_JTLA3 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLA3 = 2.0678e-15
.param B0_JTLA3 = 1
.param Ic0_JTLA3 = 1.0000e-04
.param IcRs_JTLA3 = 6.8599e-04
.param B0Rs_JTLA3 = 6.8599
.param Rsheet_JTLA3 = 2
.param Lsheet_JTLA3 = 1.1300e-12
.param LP_JTLA3 = 2.0000e-13
.param IC_JTLA3 = 2.5000
.param Lptl_JTLA3 = 2.0000e-12
.param LB_JTLA3 = 2.0000e-12
.param BiasCoef_JTLA3 = 0.7000
.param B1_JTLA3 = 2.5000
.param B2_JTLA3 = 2.5000
.param IB1_JTLA3 = 3.5000e-04
.param LB1_JTLA3 = 2.0000e-12
.param L1_JTLA3 = 2.0678e-12
.param L2_JTLA3 = 2.0678e-12
.param L3_JTLA3 = 2.0678e-12
.param L4_JTLA3 = 2.0678e-12
.param RB1_JTLA3 = 2.7440
.param RB2_JTLA3 = 2.7440
.param LRB1_JTLA3 = 1.7503e-12
.param LRB2_JTLA3 = 1.7503e-12
.param LP1_JTLA3 = 2.0000e-13
.param LP2_JTLA3 = 2.0000e-13

B1_JTLA3 1_JTLA3 2_JTLA3 jjmit_JTLA3 area=B1_JTLA3
B2_JTLA3 6_JTLA3 7_JTLA3 jjmit_JTLA3 area=B2_JTLA3
IB1_JTLA3 0 5_JTLA3 pwl(0 0 5p IB1_JTLA3)
L1_JTLA3 a_JTLA3 1_JTLA3 2.082E-12
L2_JTLA3 1_JTLA3 4_JTLA3 2.06E-12
L3_JTLA3 4_JTLA3 6_JTLA3 2.067E-12
L4_JTLA3 6_JTLA3 q_JTLA3 2.075E-12
LP1_JTLA3 2_JTLA3 0 4.998E-13
LP2_JTLA3 7_JTLA3 0 5.011E-13
LB1_JTLA3 5_JTLA3 4_JTLA3 LB1_JTLA3
RB1_JTLA3 1_JTLA3 3_JTLA3 RB1_JTLA3
RB2_JTLA3 6_JTLA3 8_JTLA3 RB2_JTLA3
LRB1_JTLA3 3_JTLA3 0 LRB1_JTLA3
LRB2_JTLA3 8_JTLA3 0 LRB2_JTLA3

*JTLA4
LC_JTLA4_1 OR2 a_JTLA4 0
LC_JTLA4_2 OR3 q_JTLA4 0

.model jjmit_JTLA4 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTLA4 = 2.0678e-15
.param B0_JTLA4 = 1
.param Ic0_JTLA4 = 1.0000e-04
.param IcRs_JTLA4 = 6.8599e-04
.param B0Rs_JTLA4 = 6.8599
.param Rsheet_JTLA4 = 2
.param Lsheet_JTLA4 = 1.1300e-12
.param LP_JTLA4 = 2.0000e-13
.param IC_JTLA4 = 2.5000
.param Lptl_JTLA4 = 2.0000e-12
.param LB_JTLA4 = 2.0000e-12
.param BiasCoef_JTLA4 = 0.7000
.param B1_JTLA4 = 2.5000
.param B2_JTLA4 = 2.5000
.param IB1_JTLA4 = 3.5000e-04
.param LB1_JTLA4 = 2.0000e-12
.param L1_JTLA4 = 2.0678e-12
.param L2_JTLA4 = 2.0678e-12
.param L3_JTLA4 = 2.0678e-12
.param L4_JTLA4 = 2.0678e-12
.param RB1_JTLA4 = 2.7440
.param RB2_JTLA4 = 2.7440
.param LRB1_JTLA4 = 1.7503e-12
.param LRB2_JTLA4 = 1.7503e-12
.param LP1_JTLA4 = 2.0000e-13
.param LP2_JTLA4 = 2.0000e-13

B1_JTLA4 1_JTLA4 2_JTLA4 jjmit_JTLA4 area=B1_JTLA4
B2_JTLA4 6_JTLA4 7_JTLA4 jjmit_JTLA4 area=B2_JTLA4
IB1_JTLA4 0 5_JTLA4 pwl(0 0 5p IB1_JTLA4)
L1_JTLA4 a_JTLA4 1_JTLA4 2.082E-12
L2_JTLA4 1_JTLA4 4_JTLA4 2.06E-12
L3_JTLA4 4_JTLA4 6_JTLA4 2.067E-12
L4_JTLA4 6_JTLA4 q_JTLA4 2.075E-12
LP1_JTLA4 2_JTLA4 0 4.998E-13
LP2_JTLA4 7_JTLA4 0 5.011E-13
LB1_JTLA4 5_JTLA4 4_JTLA4 LB1_JTLA4
RB1_JTLA4 1_JTLA4 3_JTLA4 RB1_JTLA4
RB2_JTLA4 6_JTLA4 8_JTLA4 RB2_JTLA4
LRB1_JTLA4 3_JTLA4 0 LRB1_JTLA4
LRB2_JTLA4 8_JTLA4 0 LRB2_JTLA4




*AND1

LC_and1_1 A1 a_and1 0
LC_and1_2 B1 b_and1 0
LC_and1_3 AND1 Q_and1 0

.param b1_and1 = 1.39878486e+00
.param bd1_and1 = 1.38855937e+00
.param l1_and1 = 1.64204687e-12
.param rd1_and1 = 6.00718616e-01
.param i1_and1 = 1.54457273e-05
.param b3_and1 = 1.51517089e+00
*This line was edited to make the simulation work
*This might change the whole margins of the file. Need to check if AND is still okay with this.
.param l3_and1 = 4.24567618e-13
.param rh1_and1 = 4.76237371e+00
.param ldp1_and1 = 1e-12
.param b2_and1 = b1_and1
.param bd2_and1 = bd1_and1
.param l2_and1 = l1_and1
.param ldp2_and1 = ldp1_and1
.param rd2_and1 = rd1_and1
.param lp1_and1 = 0.2e-12
.param lhp1_and1 = 1e-12
.param lhp2_and1 = lhp1_and1
.param rh2_and1 = rh1_and1

.model jjmit_and1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

b1_and1 30_and1 10_and1 jjmit_and1 area=b1_and1
b2_and1 30_and1 20_and1 jjmit_and1 area=b2_and1
b3_and1 31_and1 30_and1 jjmit_and1 area=b3_and1
bd1_and1 30_and1 12_and1 jjmit_and1 area=bd1_and1
bd2_and1 30_and1 22_and1 jjmit_and1 area=bd2_and1
i1_and1 0 30_and1 pwl(0 0 5p i1_and1)
l1_and1 A_and1 10_and1 l1_and1
l2_and1 B_and1 20_and1 l2_and1
l3_and1 30_and1 Q_and1 l3_and1
ldp1_and1 11_and1 12_and1 ldp1_and1
ldp2_and1 21_and1 22_and1 ldp2_and1
lhp1_and1 13_and1 30_and1 lhp1_and1
lhp2_and1 23_and1 30_and1 lhp2_and1
lp1_and1 31_and1 0 lp1_and1
rd1_and1 11_and1 10_and1 rd1_and1
rd2_and1 21_and1 20_and1 rd2_and1
rh1_and1 13_and1 10_and1 rh1_and1
rh2_and1 23_and1 20_and1 rh2_and1


*AND2

LC_and2_1 AND2 a_and2 0
LC_and2_2 OR3 b_and2 0
LC_and2_3 Q Q_and2 0

.param b1_and2 = 1.39878486e+00
.param bd1_and2 = 1.38855937e+00
.param l1_and2 = 1.64204687e-12
.param rd1_and2 = 6.00718616e-01
.param i1_and2 = 1.54457273e-05
.param b3_and2 = 1.51517089e+00
*This line was edited to make the simulation work
*This might change the whole margins of the file. Need to check if AND is still okay with this.
.param l3_and2 = 4.24567618e-13
.param rh1_and2 = 4.76237371e+00
.param ldp1_and2 = 1e-12
.param b2_and2 = b1_and2
.param bd2_and2 = bd1_and2
.param l2_and2 = l1_and2
.param ldp2_and2 = ldp1_and2
.param rd2_and2 = rd1_and2
.param lp1_and2 = 0.2e-12
.param lhp1_and2 = 1e-12
.param lhp2_and2 = lhp1_and2
.param rh2_and2 = rh1_and2

.model jjmit_and2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)

b1_and2 30_and2 10_and2 jjmit_and2 area=b1_and2
b2_and2 30_and2 20_and2 jjmit_and2 area=b2_and2
b3_and2 31_and2 30_and2 jjmit_and2 area=b3_and2
bd1_and2 30_and2 12_and2 jjmit_and2 area=bd1_and2
bd2_and2 30_and2 22_and2 jjmit_and2 area=bd2_and2
i1_and2 0 30_and2 pwl(0 0 5p i1_and2)
l1_and2 A_and2 10_and2 l1_and2
l2_and2 B_and2 20_and2 l2_and2
l3_and2 30_and2 Q_and2 l3_and2
ldp1_and2 11_and2 12_and2 ldp1_and2
ldp2_and2 21_and2 22_and2 ldp2_and2
lhp1_and2 13_and2 30_and2 lhp1_and2
lhp2_and2 23_and2 30_and2 lhp2_and2
lp1_and2 31_and2 0 lp1_and2
rd1_and2 11_and2 10_and2 rd1_and2
rd2_and2 21_and2 20_and2 rd2_and2
rh1_and2 13_and2 10_and2 rh1_and2
rh2_and2 23_and2 20_and2 rh2_and2




* XOR     DSFQ_ORi     A1     B2   OR1

LC_OR1_1 A1 a_OR1 0
LC_OR1_2 B2 b_OR1 0
LC_OR1_3 OR1 Q_OR1 0

* .subckt DSFQ_OR1 a_OR1 b_OR1 q_OR1
.model jjmit_OR1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
*Confluence Buffer A
.param l1_OR1 = 2e-12
.param b1_OR1 = 1.37211310e+00
.param b3_OR1 = 2.77209629e+00
.param b4_OR1 = 3.78734058e-01

* AND GATE LOOP
.param l4_OR1 = 1.22182342e-12
.param b7_OR1 = 1.19265113e+00
.param b9_OR1 = 5.40924075e-01
.param l7_OR1 = 1.62539785e-13
.param r1_OR1 = 1.09745275e+01
.param r2_OR1 = 5.58089917e-01
.param l5_OR1 = 5.61756493e-13

* Output Stage
.param b8_OR1 = 7.09413113e-01
.param i1_OR1 = 3.23631555e-04
.param l3_OR1 = 2e-12
.param l6_OR1 = 3.06315548e-12

*Confluence Buffer B
.param l2_OR1 = L1_OR1
.param b2_OR1 = B1_OR1
.param b5_OR1 = B3_OR1
.param b6_OR1 = B4_OR1

*Parasitics
.param lp1_OR1 = 0.2e-12
.param lp2_OR1 = 0.2e-12
.param lp3_OR1 = 0.2e-12
.param lp4_OR1 = 0.2e-12

* Back Annotated .cir file from KiCad
b1_OR1 3_OR1 1_OR1 jjmit_OR1 area=b1_OR1
b2_OR1 4_OR1 2_OR1 jjmit_OR1 area=b2_OR1
b3_OR1 3_OR1 10_OR1 jjmit_OR1 area=b3_OR1
b4_OR1 5_OR1 3_OR1 jjmit_OR1 area=b4_OR1
b5_OR1 4_OR1 10_OR1 jjmit_OR1 area=b5_OR1
b6_OR1 6_OR1 4_OR1 jjmit_OR1 area=b6_OR1
b7_OR1 24_OR1 20_OR1 jjmit_OR1 area=b7_OR1
b8_OR1 30_OR1 31_OR1 jjmit_OR1 area=b8_OR1
b9_OR1 24_OR1 23_OR1 jjmit_OR1 area=b9_OR1
i1_OR1 0 10_OR1 pwl(0 0 5p i1_OR1)
l1_OR1 a_OR1 1_OR1 l1_OR1
l2_OR1 b_OR1 2_OR1 l2_OR1
l3_OR1 10_OR1 30_OR1 l3_OR1
l4_OR1 30_OR1 20_OR1 l4_OR1
l5_OR1 21_OR1 24_OR1 l5_OR1
l6_OR1 30_OR1 q_OR1 l6_OR1
l7_OR1 22_OR1 23_OR1 l7_OR1
lp1_OR1 5_OR1 0 lp1_OR1
lp2_OR1 6_OR1 0 lp2_OR1
lp3_OR1 24_OR1 0 lp3_OR1
lp4_OR1 31_OR1 0 lp4_OR1
r1_OR1 21_OR1 20_OR1 r1_OR1
r2_OR1 22_OR1 20_OR1 r2_OR1




* XNAND2  DSFQ_NOTo    AND1   A11   B11   AND2

LC_NOT_1 Annn AND1 0
LC_NOT_2 Bnnn A11 0
LC_NOT_3 Cnnn B11 0
LC_NOT_4 Qnnn AND2 0

*************** NEW NOT GATE
* .subckt DSFQ_NOTo A B C Q
* .model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
*A is inverting input.
*B and C are inputs for the OR gate.
*Q is output.

* XDSFQ_OR DSFQ_ORi B C CLKD
* XJTLCLK LSMITLL_JTLi CLKD CLK
* XNOTLS LSMITLL_NOTi A CLK Q

*NNOT

LC_NOT_NOT_1 Annn a_NOT_NOT 0
LC_NOT_NOT_2 CLK clk_NOT_NOT 0
LC_NOT_NOT_3 Qnnn q_NOT_NOT 0
* .subckt LSMITLL_NOTi_NOT_NOT a_NOT_NOT clk_NOT_NOT q_NOT_NOT
.model jjmit_NOT_NOT jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_NOT_NOT = 2.0678e-15
.param B0_NOT_NOT = 1
.param Ic0_NOT_NOT = 1.0000e-04
.param IcRs_NOT_NOT = 6.8599e-04
.param B0Rs_NOT_NOT = 6.8599
.param Rsheet_NOT_NOT = 2
.param Lsheet_NOT_NOT = 1.1300e-12
.param LP_NOT_NOT = 2.0000e-13
.param IC_NOT_NOT = 2.5000
.param LB_NOT_NOT = 2.0000e-12
.param BiasCoef_NOT_NOT = 0.7000
.param B1_NOT_NOT = 2.5000
.param B2_NOT_NOT = 2.5700
.param B3_NOT_NOT = 1.0700
.param B4_NOT_NOT = 2.5000
.param B5_NOT_NOT = 1.3400
.param B6_NOT_NOT = 3.0300
.param B7_NOT_NOT = 1.3800
.param B8_NOT_NOT = 0.8000
.param B9_NOT_NOT = 2.5000
.param IB1_NOT_NOT = 1.7500e-04
.param IB2_NOT_NOT = 8.7000e-05
.param IB3_NOT_NOT = 2.5700e-04
.param IB4_NOT_NOT = 1.7500e-04
.param IB5_NOT_NOT = 1.7500e-04
.param LB1_NOT_NOT = 2.0000e-12
.param LB2_NOT_NOT = 2.0000e-12
.param LB3_NOT_NOT = 2.0000e-12
.param LB4_NOT_NOT = 2.0000e-12
.param LB5_NOT_NOT = 2.0000e-12
.param RB1_NOT_NOT = 2.7440
.param RB2_NOT_NOT = 2.6692
.param RB3_NOT_NOT = 6.4111
.param RB4_NOT_NOT = 2.7440
.param RB5_NOT_NOT = 5.1193
.param RB6_NOT_NOT = 2.2640
.param RB7_NOT_NOT = 4.9709
.param RB8_NOT_NOT = 8.5749
.param RB9_NOT_NOT = 2.7440
.param LRB1_NOT_NOT = 1.5503e-12
.param LRB2_NOT_NOT = 1.5081e-12
.param LRB3_NOT_NOT = 3.6223e-12
.param LRB4_NOT_NOT = 1.5503e-12
.param LRB5_NOT_NOT = 2.8924e-12
.param LRB6_NOT_NOT = 1.2792e-12
.param LRB7_NOT_NOT = 2.8086e-12
.param LRB8_NOT_NOT = 4.8448e-12
.param LRB9_NOT_NOT = 1.5503e-12
.param RD_NOT_NOT = 4
.param LRD_NOT_NOT = 2.0000e-12

B1_NOT_NOT 1_NOT_NOT 2_NOT_NOT jjmit_NOT_NOT area=B1_NOT_NOT
B2_NOT_NOT 4_NOT_NOT 5_NOT_NOT jjmit_NOT_NOT area=B2_NOT_NOT
B3_NOT_NOT 7_NOT_NOT 8_NOT_NOT jjmit_NOT_NOT area=B3_NOT_NOT
B4_NOT_NOT 13_NOT_NOT 14_NOT_NOT jjmit_NOT_NOT area=B4_NOT_NOT
B5_NOT_NOT 17_NOT_NOT 18_NOT_NOT jjmit_NOT_NOT area=B5_NOT_NOT
B6_NOT_NOT 10_NOT_NOT 11_NOT_NOT jjmit_NOT_NOT area=B6_NOT_NOT
B7_NOT_NOT 20_NOT_NOT 18_NOT_NOT jjmit_NOT_NOT area=B7_NOT_NOT
B8_NOT_NOT 18_NOT_NOT 19_NOT_NOT jjmit_NOT_NOT area=B8_NOT_NOT
B9_NOT_NOT 21_NOT_NOT 22_NOT_NOT jjmit_NOT_NOT area=B9_NOT_NOT

IB1_NOT_NOT 0 3_NOT_NOT pwl(0 0 5p IB1_NOT_NOT)
IB2_NOT_NOT 0 6_NOT_NOT pwl(0 0 5p IB2_NOT_NOT)
IB3_NOT_NOT 0 9_NOT_NOT pwl(0 0 5p IB3_NOT_NOT)
IB4_NOT_NOT 0 15_NOT_NOT pwl(0 0 5p IB4_NOT_NOT)
IB5_NOT_NOT 0 23_NOT_NOT pwl(0 0 5p IB5_NOT_NOT)

LB1_NOT_NOT 3_NOT_NOT 1_NOT_NOT LB1_NOT_NOT
LB2_NOT_NOT 6_NOT_NOT 4_NOT_NOT LB2_NOT_NOT
LB3_NOT_NOT 8_NOT_NOT 9_NOT_NOT LB3_NOT_NOT
LB4_NOT_NOT 13_NOT_NOT 15_NOT_NOT LB4_NOT_NOT
LB5_NOT_NOT 21_NOT_NOT 23_NOT_NOT LB5_NOT_NOT

L1_NOT_NOT a_NOT_NOT 1_NOT_NOT 2.062E-12
L2_NOT_NOT 1_NOT_NOT 4_NOT_NOT 1.889E-12
L3_NOT_NOT 4_NOT_NOT 7_NOT_NOT 2.72E-12
L4_NOT_NOT clk_NOT_NOT 13_NOT_NOT 2.057E-12
L5_NOT_NOT 13_NOT_NOT 16_NOT_NOT 1.029E-12
L6_NOT_NOT 16_NOT_NOT 17_NOT_NOT 1.241E-12
L7_NOT_NOT 16_NOT_NOT 12_NOT_NOT 1.973E-12
L8_NOT_NOT 10_NOT_NOT 12_NOT_NOT 1.003E-12
L9_NOT_NOT 10_NOT_NOT 8_NOT_NOT 7.524E-12
L10_NOT_NOT 8_NOT_NOT 20_NOT_NOT 1.234E-12
L11_NOT_NOT 18_NOT_NOT 21_NOT_NOT 2.607E-12
L12_NOT_NOT 21_NOT_NOT q_NOT_NOT 2.062E-12

LP1_NOT_NOT 2_NOT_NOT 0 5.271E-13
LP2_NOT_NOT 5_NOT_NOT 0 5.237E-13
LP4_NOT_NOT 14_NOT_NOT 0 4.759E-13
LP6_NOT_NOT 11_NOT_NOT 0 5.021E-13
LP8_NOT_NOT 19_NOT_NOT 0 6.33E-13
LP9_NOT_NOT 22_NOT_NOT 0 4.749E-13

RB1_NOT_NOT 1_NOT_NOT 101_NOT_NOT RB1_NOT_NOT
LRB1_NOT_NOT 101_NOT_NOT 0 LRB1_NOT_NOT
RB2_NOT_NOT 4_NOT_NOT 104_NOT_NOT RB2_NOT_NOT
LRB2_NOT_NOT 104_NOT_NOT 5_NOT_NOT LRB2_NOT_NOT
RB3_NOT_NOT 7_NOT_NOT 107_NOT_NOT RB3_NOT_NOT
LRB3_NOT_NOT 107_NOT_NOT 8_NOT_NOT LRB3_NOT_NOT
RB4_NOT_NOT 13_NOT_NOT 113_NOT_NOT RB4_NOT_NOT
LRB4_NOT_NOT 113_NOT_NOT 0 LRB4_NOT_NOT
RB5_NOT_NOT 17_NOT_NOT 117_NOT_NOT RB5_NOT_NOT
LRB5_NOT_NOT 117_NOT_NOT 18_NOT_NOT LRB5_NOT_NOT
RB6_NOT_NOT 10_NOT_NOT 110_NOT_NOT RB6_NOT_NOT
LRB6_NOT_NOT 110_NOT_NOT 0 LRB6_NOT_NOT
RB7_NOT_NOT 20_NOT_NOT 120_NOT_NOT RB7_NOT_NOT
LRB7_NOT_NOT 120_NOT_NOT 18_NOT_NOT LRB7_NOT_NOT
RB8_NOT_NOT 18_NOT_NOT 118_NOT_NOT RB8_NOT_NOT
LRB8_NOT_NOT 118_NOT_NOT 0 LRB8_NOT_NOT
RB9_NOT_NOT 21_NOT_NOT 121_NOT_NOT RB9_NOT_NOT
LRB9_NOT_NOT 121_NOT_NOT 0 LRB9_NOT_NOT
LRD_NOT_NOT 12_NOT_NOT 112_NOT_NOT LRD_NOT_NOT
RD_NOT_NOT 112_NOT_NOT 0 RD_NOT_NOT




*JTL_NOT

LC_JTL_NOT_1 CLKD a_JTL_NOT 0
LC_JTL_NOT_2 CLK q_JTL_NOT 0

.model jjmit_JTL_NOT jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_JTL_NOT = 2.0678e-15
.param B0_JTL_NOT = 1
.param Ic0_JTL_NOT = 1.0000e-04
.param IcRs_JTL_NOT = 6.8599e-04
.param B0Rs_JTL_NOT = 6.8599
.param Rsheet_JTL_NOT = 2
.param Lsheet_JTL_NOT = 1.1300e-12
.param LP_JTL_NOT = 2.0000e-13
.param IC_JTL_NOT = 2.5000
.param Lptl_JTL_NOT = 2.0000e-12
.param LB_JTL_NOT = 2.0000e-12
.param BiasCoef_JTL_NOT = 0.7000
.param B1_JTL_NOT = 2.5000
.param B2_JTL_NOT = 2.5000
.param IB1_JTL_NOT = 3.5000e-04
.param LB1_JTL_NOT = 2.0000e-12
.param L1_JTL_NOT = 2.0678e-12
.param L2_JTL_NOT = 2.0678e-12
.param L3_JTL_NOT = 2.0678e-12
.param L4_JTL_NOT = 2.0678e-12
.param RB1_JTL_NOT = 2.7440
.param RB2_JTL_NOT = 2.7440
.param LRB1_JTL_NOT = 1.7503e-12
.param LRB2_JTL_NOT = 1.7503e-12
.param LP1_JTL_NOT = 2.0000e-13
.param LP2_JTL_NOT = 2.0000e-13

B1_JTL_NOT 1_JTL_NOT 2_JTL_NOT jjmit_JTL_NOT area=B1_JTL_NOT
B2_JTL_NOT 6_JTL_NOT 7_JTL_NOT jjmit_JTL_NOT area=B2_JTL_NOT
IB1_JTL_NOT 0 5_JTL_NOT pwl(0 0 5p IB1_JTL_NOT)
L1_JTL_NOT a_JTL_NOT 1_JTL_NOT 2.082E-12
L2_JTL_NOT 1_JTL_NOT 4_JTL_NOT 2.06E-12
L3_JTL_NOT 4_JTL_NOT 6_JTL_NOT 2.067E-12
L4_JTL_NOT 6_JTL_NOT q_JTL_NOT 2.075E-12
LP1_JTL_NOT 2_JTL_NOT 0 4.998E-13
LP2_JTL_NOT 7_JTL_NOT 0 5.011E-13
LB1_JTL_NOT 5_JTL_NOT 4_JTL_NOT LB1_JTL_NOT
RB1_JTL_NOT 1_JTL_NOT 3_JTL_NOT RB1_JTL_NOT
RB2_JTL_NOT 6_JTL_NOT 8_JTL_NOT RB2_JTL_NOT
LRB1_JTL_NOT 3_JTL_NOT 0 LRB1_JTL_NOT
LRB2_JTL_NOT 8_JTL_NOT 0 LRB2_JTL_NOT


*OR_NOT

LC_OR_NOT_1 Bnnn a_OR_NOT 0
LC_OR_NOT_2 Cnnn b_OR_NOT 0
LC_OR_NOT_3 CLKD Q_OR_NOT 0

* .subckt DSFQ_OR_NOT a_OR_NOT b_OR_NOT q_OR_NOT
.model jjmit_OR_NOT jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
*Confluence Buffer A
.param l1_OR_NOT = 2e-12
.param b1_OR_NOT = 1.37211310e+00
.param b3_OR_NOT = 2.77209629e+00
.param b4_OR_NOT = 3.78734058e-01

* AND GATE LOOP
.param l4_OR_NOT = 1.22182342e-12
.param b7_OR_NOT = 1.19265113e+00
.param b9_OR_NOT = 5.40924075e-01
.param l7_OR_NOT = 1.62539785e-13
.param r1_OR_NOT = 1.09745275e+01
.param r2_OR_NOT = 5.58089917e-01
.param l5_OR_NOT = 5.61756493e-13

* Output Stage
.param b8_OR_NOT = 7.09413113e-01
.param i1_OR_NOT = 3.23631555e-04
.param l3_OR_NOT = 2e-12
.param l6_OR_NOT = 3.06315548e-12

*Confluence Buffer B
.param l2_OR_NOT = L1_OR_NOT
.param b2_OR_NOT = B1_OR_NOT
.param b5_OR_NOT = B3_OR_NOT
.param b6_OR_NOT = B4_OR_NOT

*Parasitics
.param lp1_OR_NOT = 0.2e-12
.param lp2_OR_NOT = 0.2e-12
.param lp3_OR_NOT = 0.2e-12
.param lp4_OR_NOT = 0.2e-12

* Back Annotated .cir file from KiCad
b1_OR_NOT 3_OR_NOT 1_OR_NOT jjmit_OR_NOT area=b1_OR_NOT
b2_OR_NOT 4_OR_NOT 2_OR_NOT jjmit_OR_NOT area=b2_OR_NOT
b3_OR_NOT 3_OR_NOT 10_OR_NOT jjmit_OR_NOT area=b3_OR_NOT
b4_OR_NOT 5_OR_NOT 3_OR_NOT jjmit_OR_NOT area=b4_OR_NOT
b5_OR_NOT 4_OR_NOT 10_OR_NOT jjmit_OR_NOT area=b5_OR_NOT
b6_OR_NOT 6_OR_NOT 4_OR_NOT jjmit_OR_NOT area=b6_OR_NOT
b7_OR_NOT 24_OR_NOT 20_OR_NOT jjmit_OR_NOT area=b7_OR_NOT
b8_OR_NOT 30_OR_NOT 31_OR_NOT jjmit_OR_NOT area=b8_OR_NOT
b9_OR_NOT 24_OR_NOT 23_OR_NOT jjmit_OR_NOT area=b9_OR_NOT
i1_OR_NOT 0 10_OR_NOT pwl(0 0 5p i1_OR_NOT)
l1_OR_NOT a_OR_NOT 1_OR_NOT l1_OR_NOT
l2_OR_NOT b_OR_NOT 2_OR_NOT l2_OR_NOT
l3_OR_NOT 10_OR_NOT 30_OR_NOT l3_OR_NOT
l4_OR_NOT 30_OR_NOT 20_OR_NOT l4_OR_NOT
l5_OR_NOT 21_OR_NOT 24_OR_NOT l5_OR_NOT
l6_OR_NOT 30_OR_NOT q_OR_NOT l6_OR_NOT
l7_OR_NOT 22_OR_NOT 23_OR_NOT l7_OR_NOT
lp1_OR_NOT 5_OR_NOT 0 lp1_OR_NOT
lp2_OR_NOT 6_OR_NOT 0 lp2_OR_NOT
lp3_OR_NOT 24_OR_NOT 0 lp3_OR_NOT
lp4_OR_NOT 31_OR_NOT 0 lp4_OR_NOT
r1_OR_NOT 21_OR_NOT 20_OR_NOT r1_OR_NOT
r2_OR_NOT 22_OR_NOT 20_OR_NOT r2_OR_NOT


*** SPLIT CELLS********************************************************************************************************************************

LC_split1_1 A a_split1 0
LC_split1_2 A1 q0_split1 0
LC_split1_3 A2 q1_split1 0
.model jjmit_split1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_split1 = 2.0678e-15
.param B0_split1 = 1
.param Ic0_split1 = 1.0000e-04
.param IcRs_split1 = 6.8599e-04
.param B0Rs_split1 = 6.8599
.param Rsheet_split1 = 2
.param Lsheet_split1 = 1.1300e-12
.param LP_split1 = 2.0000e-13
.param IC_split1 = 2.5000
.param Lptl_split1 = 2.0000e-12
.param LB_split1 = 2.0000e-12
.param BiasCoef_split1 = 0.7000
.param RD_split1 = 1.3600
.param B1_split1 = 2.5000
.param B2_split1 = 3
.param B3_split1 = 2.5000
.param B4_split1 = 2.5000
.param IB1_split1 = 1.7500e-04
.param IB2_split1 = 2.8000e-04
.param IB3_split1 = 1.7500e-04
.param IB4_split1 = 1.7500e-04
.param L1_split1 = 2.0000e-12
.param L2_split1 = 4.1357e-12
.param L3_split1 = 1.7232e-12
.param L4_split1 = 1.7232e-12
.param L5_split1 = 2.0000e-12
.param L6_split1 = 1.7232e-12
.param L7_split1 = 2.0000e-12
.param RB1_split1 = 2.7440
.param RB2_split1 = 2.2866
.param RB3_split1 = 2.7440
.param RB4_split1 = 2.7440
.param LRB1_split1 = 1.5503e-12
.param LRB2_split1 = 1.2919e-12
.param LRB3_split1 = 1.5503e-12
.param LRB4_split1 = 1.5503e-12

IB1_split1 0 3_split1 pwl(0 0 5p IB1_split1)
IB2_split1 0 6_split1 pwl(0 0 5p IB2_split1)
IB3_split1 0 10_split1 pwl(0 0 5p IB3_split1)
IB4_split1 0 13_split1 pwl(0 0 5p IB4_split1)
LB1_split1 3_split1 1_split1 9.175E-13
LB2_split1 6_split1 4_split1 7.666E-13
LB3_split1 10_split1 8_split1 1.928E-12
LB4_split1 13_split1 11_split1 8.786E-13

B1_split1 1_split1 2_split1 jjmit_split1 area=B1_split1
B2_split1 4_split1 5_split1 jjmit_split1 area=B2_split1
B3_split1 8_split1 9_split1 jjmit_split1 area=B3_split1
B4_split1 11_split1 12_split1 jjmit_split1 area=B4_split1
L1_split1 a_split1 1_split1 2.063E-12
L2_split1 1_split1 4_split1 3.637E-12
L3_split1 4_split1 7_split1 1.278E-12
L4_split1 7_split1 8_split1 1.305E-12
L5_split1 8_split1 q0_split1 2.05E-12
L6_split1 7_split1 11_split1 1.315E-12
L7_split1 11_split1 q1_split1 2.06E-12

LP1_split1 2_split1 0 4.676E-13
LP2_split1 5_split1 0 4.498E-13
LP3_split1 9_split1 0 5.183E-13
LP4_split1 12_split1 0 4.639E-13
RB1_split1 1_split1 101_split1 RB1_split1
LRB1_split1 101_split1 0 LRB1_split1
RB2_split1 4_split1 104_split1 RB2_split1
LRB2_split1 104_split1 0 LRB2_split1
RB3_split1 8_split1 108_split1 RB3_split1
LRB3_split1 108_split1 0 LRB3_split1
RB4_split1 11_split1 111_split1 RB4_split1
LRB4_split1 111_split1 0 LRB4_split1



*SPLIT2



LC_split2_1 B a_split2 0
LC_split2_2 B1 q0_split2 0
LC_split2_3 B2 q1_split2 0
.model jjmit_split2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0_split2 = 2.0678e-15
.param B0_split2 = 1
.param Ic0_split2 = 1.0000e-04
.param IcRs_split2 = 6.8599e-04
.param B0Rs_split2 = 6.8599
.param Rsheet_split2 = 2
.param Lsheet_split2 = 1.1300e-12
.param LP_split2 = 2.0000e-13
.param IC_split2 = 2.5000
.param Lptl_split2 = 2.0000e-12
.param LB_split2 = 2.0000e-12
.param BiasCoef_split2 = 0.7000
.param RD_split2 = 1.3600
.param B1_split2 = 2.5000
.param B2_split2 = 3
.param B3_split2 = 2.5000
.param B4_split2 = 2.5000
.param IB1_split2 = 1.7500e-04
.param IB2_split2 = 2.8000e-04
.param IB3_split2 = 1.7500e-04
.param IB4_split2 = 1.7500e-04
.param L1_split2 = 2.0000e-12
.param L2_split2 = 4.1357e-12
.param L3_split2 = 1.7232e-12
.param L4_split2 = 1.7232e-12
.param L5_split2 = 2.0000e-12
.param L6_split2 = 1.7232e-12
.param L7_split2 = 2.0000e-12
.param RB1_split2 = 2.7440
.param RB2_split2 = 2.2866
.param RB3_split2 = 2.7440
.param RB4_split2 = 2.7440
.param LRB1_split2 = 1.5503e-12
.param LRB2_split2 = 1.2919e-12
.param LRB3_split2 = 1.5503e-12
.param LRB4_split2 = 1.5503e-12

IB1_split2 0 3_split2 pwl(0 0 5p IB1_split2)
IB2_split2 0 6_split2 pwl(0 0 5p IB2_split2)
IB3_split2 0 10_split2 pwl(0 0 5p IB3_split2)
IB4_split2 0 13_split2 pwl(0 0 5p IB4_split2)
LB1_split2 3_split2 1_split2 9.175E-13
LB2_split2 6_split2 4_split2 7.666E-13
LB3_split2 10_split2 8_split2 1.928E-12
LB4_split2 13_split2 11_split2 8.786E-13

B1_split2 1_split2 2_split2 jjmit_split2 area=B1_split2
B2_split2 4_split2 5_split2 jjmit_split2 area=B2_split2
B3_split2 8_split2 9_split2 jjmit_split2 area=B3_split2
B4_split2 11_split2 12_split2 jjmit_split2 area=B4_split2
L1_split2 a_split2 1_split2 2.063E-12
L2_split2 1_split2 4_split2 3.637E-12
L3_split2 4_split2 7_split2 1.278E-12
L4_split2 7_split2 8_split2 1.305E-12
L5_split2 8_split2 q0_split2 2.05E-12
L6_split2 7_split2 11_split2 1.315E-12
L7_split2 11_split2 q1_split2 2.06E-12

LP1_split2 2_split2 0 4.676E-13
LP2_split2 5_split2 0 4.498E-13
LP3_split2 9_split2 0 5.183E-13
LP4_split2 12_split2 0 4.639E-13
RB1_split2 1_split2 101_split2 RB1_split2
LRB1_split2 101_split2 0 LRB1_split2
RB2_split2 4_split2 104_split2 RB2_split2
LRB2_split2 104_split2 0 LRB2_split2
RB3_split2 8_split2 108_split2 RB3_split2
LRB3_split2 108_split2 0 LRB3_split2
RB4_split2 11_split2 111_split2 RB4_split2
LRB4_split2 111_split2 0 LRB4_split2

.ends